// Verilog netlist created by Tang Dynasty v5.6.119222
// Sat Oct 19 17:02:28 2024

`timescale 1ns / 1ps
module Divider_32
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [31:0] denominator;
  input [31:0] numerator;
  input rst;
  input start;
  output done;
  output [31:0] quotient;
  output [31:0] remainder;

  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 32;
  parameter W_NUM = 32;
  // localparam W_CNT = 6;
  wire [5:0] al_1deac949;
  wire [5:0] al_d0dc52fd;
  wire [5:0] al_537e4616;
  wire [62:0] al_11033702;
  wire [62:0] al_1c1b24e7;
  wire [31:0] al_1315ed94;
  wire [31:0] al_9bfb1470;
  wire [62:0] al_c67bebad;
  wire [31:0] al_327525b3;
  wire al_30a8497b;
  wire al_32d88032;
  wire al_6862943f;
  wire al_31eb4985;
  wire al_cd217c4a;
  wire al_a707256f;
  wire al_9673d977;
  wire al_a9fbe072;
  wire al_3973d008;
  wire al_4c40b6e5;
  wire al_d63e42fe;
  wire al_b4fc1000;
  wire al_ab829401;
  wire al_b7ca2ed;
  wire al_22a7ce9f;
  wire al_f5902502;
  wire al_b83a67b2;
  wire al_540b209;
  wire al_27e1f3bc;
  wire al_e64e5f1c;
  wire al_e761a920;
  wire al_42ead886;
  wire al_f5a327ab;
  wire al_b23e28b5;
  wire al_283f8d98;
  wire al_516747bd;
  wire al_88a2e01;
  wire al_424d2e3a;
  wire al_5d3a435a;
  wire al_4a5ad68f;
  wire al_9646e713;
  wire al_6cee34b4;
  wire al_9015d2c4;
  wire al_64efb4d0;
  wire al_2d9efd6f;
  wire al_e033469;
  wire al_52f68b55;
  wire al_6b2ca00d;
  wire al_92782c7;
  wire al_ba378049;
  wire al_abb07f01;
  wire al_3a3b377;
  wire al_f762b252;
  wire al_6c2df81c;
  wire al_81606498;
  wire al_fef7e453;
  wire al_84e7266e;
  wire al_5866a5aa;
  wire al_18356e63;
  wire al_4bbb767a;
  wire al_5b37f318;
  wire al_19d272d0;
  wire al_7a6c3f49;
  wire al_59d0e94d;
  wire al_1311ca2a;
  wire al_cc41fd76;
  wire al_9d116ec6;
  wire al_31a76718;
  wire al_728d165d;
  wire al_3c978099;
  wire al_806cd1d1;
  wire al_21e6aa37;
  wire al_d47fc616;
  wire al_a4c56fd2;
  wire al_3aecfb13;
  wire al_a04afdc3;
  wire al_c8596675;
  wire al_26fbd6b;
  wire al_98b263c2;
  wire al_973a6162;
  wire al_d21ff3d4;
  wire al_20da7cd1;
  wire al_4b6c2990;
  wire al_2a9315a6;
  wire al_b9c5d958;
  wire al_56630a35;
  wire al_a1b0b17a;
  wire al_7b07bb65;
  wire al_9df2af8f;
  wire al_df20ca5b;
  wire al_ab6a0e7;
  wire al_3f047599;
  wire al_b4d1b2a2;
  wire al_469cb985;
  wire al_ffb568cb;
  wire al_8f0bd67f;
  wire al_ee5c4865;
  wire al_c617ea0a;
  wire al_c36dd466;
  wire al_cbd8eebc;
  wire al_c8debd9c;
  wire al_73a2ed86;
  wire al_c8a237ee;
  wire al_2945efc4;
  wire al_a649c440;
  wire al_90e69cc8;
  wire al_25b33d0e;
  wire al_ea1005e8;
  wire al_128ecb61;
  wire al_fb8ac41d;
  wire al_f6cfbe3c;
  wire al_ec2ed332;
  wire al_114eba31;
  wire al_c61b4192;
  wire al_2ea6dadb;

  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b22ad72b (
    .a(al_1deac949[4]),
    .b(1'b0),
    .c(al_cd217c4a),
    .o({al_a707256f,al_537e4616[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_37642c3c (
    .a(al_1deac949[5]),
    .b(1'b0),
    .c(al_a707256f),
    .o({open_n0,al_537e4616[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_8a72a648 (
    .a(1'b0),
    .o({al_30a8497b,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a4d828f2 (
    .a(al_1deac949[0]),
    .b(1'b1),
    .c(al_30a8497b),
    .o({al_32d88032,al_537e4616[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8b186716 (
    .a(al_1deac949[1]),
    .b(1'b0),
    .c(al_32d88032),
    .o({al_6862943f,al_537e4616[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3d917c9c (
    .a(al_1deac949[2]),
    .b(1'b0),
    .c(al_6862943f),
    .o({al_31eb4985,al_537e4616[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e7664728 (
    .a(al_1deac949[3]),
    .b(1'b0),
    .c(al_31eb4985),
    .o({al_cd217c4a,al_537e4616[3]}));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_dc50342 (
    .a(al_2ea6dadb),
    .b(al_1deac949[0]),
    .c(al_1deac949[5]),
    .o(al_114eba31));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(C*~(A*~(E@D))))"),
    .INIT(32'hdcfcfcdc))
    al_f17cd423 (
    .a(al_2ea6dadb),
    .b(start),
    .c(al_537e4616[0]),
    .d(al_1deac949[0]),
    .e(al_1deac949[5]),
    .o(al_d0dc52fd[0]));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(A*~(E@D)))"),
    .INIT(32'h10303010))
    al_147e6a1b (
    .a(al_2ea6dadb),
    .b(start),
    .c(al_537e4616[1]),
    .d(al_1deac949[0]),
    .e(al_1deac949[5]),
    .o(al_d0dc52fd[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c8620855 (
    .a(start),
    .b(al_537e4616[2]),
    .o(al_d0dc52fd[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6614de08 (
    .a(start),
    .b(al_537e4616[3]),
    .o(al_d0dc52fd[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6dc5f615 (
    .a(start),
    .b(al_537e4616[4]),
    .o(al_d0dc52fd[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_79196817 (
    .a(al_1deac949[1]),
    .b(al_1deac949[2]),
    .c(al_1deac949[3]),
    .d(al_1deac949[4]),
    .o(al_2ea6dadb));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(A*~(E@D)))"),
    .INIT(32'h10303010))
    al_e3df142c (
    .a(al_2ea6dadb),
    .b(start),
    .c(al_537e4616[5]),
    .d(al_1deac949[0]),
    .e(al_1deac949[5]),
    .o(al_d0dc52fd[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_12c43e12 (
    .a(denominator[0]),
    .b(start),
    .c(al_11033702[32]),
    .o(al_1c1b24e7[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ded93226 (
    .a(denominator[1]),
    .b(start),
    .c(al_11033702[33]),
    .o(al_1c1b24e7[32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c35e0dcc (
    .a(denominator[2]),
    .b(start),
    .c(al_11033702[34]),
    .o(al_1c1b24e7[33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_362a2d70 (
    .a(denominator[3]),
    .b(start),
    .c(al_11033702[35]),
    .o(al_1c1b24e7[34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_619d59f3 (
    .a(denominator[4]),
    .b(start),
    .c(al_11033702[36]),
    .o(al_1c1b24e7[35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8b9da26a (
    .a(denominator[5]),
    .b(start),
    .c(al_11033702[37]),
    .o(al_1c1b24e7[36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_14645c1e (
    .a(denominator[6]),
    .b(start),
    .c(al_11033702[38]),
    .o(al_1c1b24e7[37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_41e73ba7 (
    .a(denominator[7]),
    .b(start),
    .c(al_11033702[39]),
    .o(al_1c1b24e7[38]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1a059b5b (
    .a(denominator[8]),
    .b(start),
    .c(al_11033702[40]),
    .o(al_1c1b24e7[39]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e68968e1 (
    .a(denominator[9]),
    .b(start),
    .c(al_11033702[41]),
    .o(al_1c1b24e7[40]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_9ae2b38c (
    .a(denominator[10]),
    .b(start),
    .c(al_11033702[42]),
    .o(al_1c1b24e7[41]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c5a5b946 (
    .a(denominator[11]),
    .b(start),
    .c(al_11033702[43]),
    .o(al_1c1b24e7[42]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7885a4da (
    .a(denominator[12]),
    .b(start),
    .c(al_11033702[44]),
    .o(al_1c1b24e7[43]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d4d1b5a8 (
    .a(denominator[13]),
    .b(start),
    .c(al_11033702[45]),
    .o(al_1c1b24e7[44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8180372b (
    .a(denominator[14]),
    .b(start),
    .c(al_11033702[46]),
    .o(al_1c1b24e7[45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f5c2596c (
    .a(denominator[15]),
    .b(start),
    .c(al_11033702[47]),
    .o(al_1c1b24e7[46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_21badd87 (
    .a(denominator[16]),
    .b(start),
    .c(al_11033702[48]),
    .o(al_1c1b24e7[47]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1f53bb72 (
    .a(denominator[17]),
    .b(start),
    .c(al_11033702[49]),
    .o(al_1c1b24e7[48]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b0febaf3 (
    .a(denominator[18]),
    .b(start),
    .c(al_11033702[50]),
    .o(al_1c1b24e7[49]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1278d55d (
    .a(denominator[19]),
    .b(start),
    .c(al_11033702[51]),
    .o(al_1c1b24e7[50]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_edab9316 (
    .a(denominator[20]),
    .b(start),
    .c(al_11033702[52]),
    .o(al_1c1b24e7[51]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1732f7be (
    .a(denominator[21]),
    .b(start),
    .c(al_11033702[53]),
    .o(al_1c1b24e7[52]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a0c3193 (
    .a(denominator[22]),
    .b(start),
    .c(al_11033702[54]),
    .o(al_1c1b24e7[53]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7ac48cbe (
    .a(denominator[23]),
    .b(start),
    .c(al_11033702[55]),
    .o(al_1c1b24e7[54]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1580b4d7 (
    .a(denominator[24]),
    .b(start),
    .c(al_11033702[56]),
    .o(al_1c1b24e7[55]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b676dfb6 (
    .a(denominator[25]),
    .b(start),
    .c(al_11033702[57]),
    .o(al_1c1b24e7[56]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a1d1fbd0 (
    .a(denominator[26]),
    .b(start),
    .c(al_11033702[58]),
    .o(al_1c1b24e7[57]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_95aaa47a (
    .a(denominator[27]),
    .b(start),
    .c(al_11033702[59]),
    .o(al_1c1b24e7[58]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1eec55a5 (
    .a(denominator[28]),
    .b(start),
    .c(al_11033702[60]),
    .o(al_1c1b24e7[59]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8c58688c (
    .a(denominator[29]),
    .b(start),
    .c(al_11033702[61]),
    .o(al_1c1b24e7[60]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_99dd0529 (
    .a(denominator[30]),
    .b(start),
    .c(al_11033702[62]),
    .o(al_1c1b24e7[61]));
  AL_DFF_0 al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_114eba31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    al_2c0796e5 (
    .a(1'b1),
    .o({al_9673d977,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c203f32c (
    .a(al_11033702[4]),
    .b(al_1315ed94[4]),
    .c(al_d63e42fe),
    .o({al_b4fc1000,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_32e253fa (
    .a(al_11033702[49]),
    .b(1'b0),
    .c(al_cc41fd76),
    .o({al_9d116ec6,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_17283bfe (
    .a(al_11033702[50]),
    .b(1'b0),
    .c(al_9d116ec6),
    .o({al_31a76718,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_99897af (
    .a(al_11033702[51]),
    .b(1'b0),
    .c(al_31a76718),
    .o({al_728d165d,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_393be1f9 (
    .a(al_11033702[52]),
    .b(1'b0),
    .c(al_728d165d),
    .o({al_3c978099,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_51bcba86 (
    .a(al_11033702[53]),
    .b(1'b0),
    .c(al_3c978099),
    .o({al_806cd1d1,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4193e874 (
    .a(al_11033702[54]),
    .b(1'b0),
    .c(al_806cd1d1),
    .o({al_21e6aa37,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3eaf5f9c (
    .a(al_11033702[55]),
    .b(1'b0),
    .c(al_21e6aa37),
    .o({al_d47fc616,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c5566d1d (
    .a(al_11033702[56]),
    .b(1'b0),
    .c(al_d47fc616),
    .o({al_a4c56fd2,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9eddbd1b (
    .a(al_11033702[57]),
    .b(1'b0),
    .c(al_a4c56fd2),
    .o({al_3aecfb13,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_245f999 (
    .a(al_11033702[58]),
    .b(1'b0),
    .c(al_3aecfb13),
    .o({al_a04afdc3,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_5a2e66a8 (
    .a(al_11033702[5]),
    .b(al_1315ed94[5]),
    .c(al_b4fc1000),
    .o({al_ab829401,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e21d4825 (
    .a(al_11033702[59]),
    .b(1'b0),
    .c(al_a04afdc3),
    .o({al_c8596675,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ef5c91b6 (
    .a(al_11033702[60]),
    .b(1'b0),
    .c(al_c8596675),
    .o({al_26fbd6b,open_n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b2778311 (
    .a(al_11033702[61]),
    .b(1'b0),
    .c(al_26fbd6b),
    .o({al_98b263c2,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ae943c46 (
    .a(al_11033702[62]),
    .b(1'b0),
    .c(al_98b263c2),
    .o({al_973a6162,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_303727b2 (
    .a(1'b0),
    .b(1'b1),
    .c(al_973a6162),
    .o({open_n23,al_c61b4192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_2f287d12 (
    .a(al_11033702[6]),
    .b(al_1315ed94[6]),
    .c(al_ab829401),
    .o({al_b7ca2ed,open_n24}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9ce86edd (
    .a(al_11033702[7]),
    .b(al_1315ed94[7]),
    .c(al_b7ca2ed),
    .o({al_22a7ce9f,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_29f6525 (
    .a(al_11033702[8]),
    .b(al_1315ed94[8]),
    .c(al_22a7ce9f),
    .o({al_f5902502,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f171b4f4 (
    .a(al_11033702[0]),
    .b(al_1315ed94[0]),
    .c(al_9673d977),
    .o({al_a9fbe072,open_n27}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e9c7012b (
    .a(al_11033702[9]),
    .b(al_1315ed94[9]),
    .c(al_f5902502),
    .o({al_b83a67b2,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4226b3d1 (
    .a(al_11033702[10]),
    .b(al_1315ed94[10]),
    .c(al_b83a67b2),
    .o({al_540b209,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3f6fc47e (
    .a(al_11033702[11]),
    .b(al_1315ed94[11]),
    .c(al_540b209),
    .o({al_27e1f3bc,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e17073e0 (
    .a(al_11033702[12]),
    .b(al_1315ed94[12]),
    .c(al_27e1f3bc),
    .o({al_e64e5f1c,open_n31}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ba5a9770 (
    .a(al_11033702[13]),
    .b(al_1315ed94[13]),
    .c(al_e64e5f1c),
    .o({al_e761a920,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cb976531 (
    .a(al_11033702[14]),
    .b(al_1315ed94[14]),
    .c(al_e761a920),
    .o({al_42ead886,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e5cd5640 (
    .a(al_11033702[15]),
    .b(al_1315ed94[15]),
    .c(al_42ead886),
    .o({al_f5a327ab,open_n34}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e4d1cd55 (
    .a(al_11033702[16]),
    .b(al_1315ed94[16]),
    .c(al_f5a327ab),
    .o({al_b23e28b5,open_n35}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_dc7e8c2c (
    .a(al_11033702[17]),
    .b(al_1315ed94[17]),
    .c(al_b23e28b5),
    .o({al_283f8d98,open_n36}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9ed345ca (
    .a(al_11033702[18]),
    .b(al_1315ed94[18]),
    .c(al_283f8d98),
    .o({al_516747bd,open_n37}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_441ad9b2 (
    .a(al_11033702[1]),
    .b(al_1315ed94[1]),
    .c(al_a9fbe072),
    .o({al_3973d008,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_36cc28eb (
    .a(al_11033702[19]),
    .b(al_1315ed94[19]),
    .c(al_516747bd),
    .o({al_88a2e01,open_n39}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e18ee10 (
    .a(al_11033702[20]),
    .b(al_1315ed94[20]),
    .c(al_88a2e01),
    .o({al_424d2e3a,open_n40}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_99bd7325 (
    .a(al_11033702[21]),
    .b(al_1315ed94[21]),
    .c(al_424d2e3a),
    .o({al_5d3a435a,open_n41}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8aa83152 (
    .a(al_11033702[22]),
    .b(al_1315ed94[22]),
    .c(al_5d3a435a),
    .o({al_4a5ad68f,open_n42}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1c94cea5 (
    .a(al_11033702[23]),
    .b(al_1315ed94[23]),
    .c(al_4a5ad68f),
    .o({al_9646e713,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_d0c6e291 (
    .a(al_11033702[24]),
    .b(al_1315ed94[24]),
    .c(al_9646e713),
    .o({al_6cee34b4,open_n44}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b1db9e6d (
    .a(al_11033702[25]),
    .b(al_1315ed94[25]),
    .c(al_6cee34b4),
    .o({al_9015d2c4,open_n45}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ada8a24f (
    .a(al_11033702[26]),
    .b(al_1315ed94[26]),
    .c(al_9015d2c4),
    .o({al_64efb4d0,open_n46}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_20b06db2 (
    .a(al_11033702[27]),
    .b(al_1315ed94[27]),
    .c(al_64efb4d0),
    .o({al_2d9efd6f,open_n47}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cbda5de1 (
    .a(al_11033702[28]),
    .b(al_1315ed94[28]),
    .c(al_2d9efd6f),
    .o({al_e033469,open_n48}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9395428b (
    .a(al_11033702[2]),
    .b(al_1315ed94[2]),
    .c(al_3973d008),
    .o({al_4c40b6e5,open_n49}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_361a841e (
    .a(al_11033702[29]),
    .b(al_1315ed94[29]),
    .c(al_e033469),
    .o({al_52f68b55,open_n50}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a4c08c3d (
    .a(al_11033702[30]),
    .b(al_1315ed94[30]),
    .c(al_52f68b55),
    .o({al_6b2ca00d,open_n51}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_d1ded6e4 (
    .a(al_11033702[31]),
    .b(al_1315ed94[31]),
    .c(al_6b2ca00d),
    .o({al_92782c7,open_n52}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f71d9d01 (
    .a(al_11033702[32]),
    .b(1'b0),
    .c(al_92782c7),
    .o({al_ba378049,open_n53}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_89b6e9ba (
    .a(al_11033702[33]),
    .b(1'b0),
    .c(al_ba378049),
    .o({al_abb07f01,open_n54}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_884478e8 (
    .a(al_11033702[34]),
    .b(1'b0),
    .c(al_abb07f01),
    .o({al_3a3b377,open_n55}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_160a5400 (
    .a(al_11033702[35]),
    .b(1'b0),
    .c(al_3a3b377),
    .o({al_f762b252,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ed8ca432 (
    .a(al_11033702[36]),
    .b(1'b0),
    .c(al_f762b252),
    .o({al_6c2df81c,open_n57}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8875c6ac (
    .a(al_11033702[37]),
    .b(1'b0),
    .c(al_6c2df81c),
    .o({al_81606498,open_n58}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3611ae8a (
    .a(al_11033702[38]),
    .b(1'b0),
    .c(al_81606498),
    .o({al_fef7e453,open_n59}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f7ac689a (
    .a(al_11033702[3]),
    .b(al_1315ed94[3]),
    .c(al_4c40b6e5),
    .o({al_d63e42fe,open_n60}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_36e3cff7 (
    .a(al_11033702[39]),
    .b(1'b0),
    .c(al_fef7e453),
    .o({al_84e7266e,open_n61}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c0e0a8b9 (
    .a(al_11033702[40]),
    .b(1'b0),
    .c(al_84e7266e),
    .o({al_5866a5aa,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1c410bbd (
    .a(al_11033702[41]),
    .b(1'b0),
    .c(al_5866a5aa),
    .o({al_18356e63,open_n63}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b713d9a8 (
    .a(al_11033702[42]),
    .b(1'b0),
    .c(al_18356e63),
    .o({al_4bbb767a,open_n64}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cf933874 (
    .a(al_11033702[43]),
    .b(1'b0),
    .c(al_4bbb767a),
    .o({al_5b37f318,open_n65}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8a1cf929 (
    .a(al_11033702[44]),
    .b(1'b0),
    .c(al_5b37f318),
    .o({al_19d272d0,open_n66}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_732efaa (
    .a(al_11033702[45]),
    .b(1'b0),
    .c(al_19d272d0),
    .o({al_7a6c3f49,open_n67}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c7d9970 (
    .a(al_11033702[46]),
    .b(1'b0),
    .c(al_7a6c3f49),
    .o({al_59d0e94d,open_n68}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a1a5dabd (
    .a(al_11033702[47]),
    .b(1'b0),
    .c(al_59d0e94d),
    .o({al_1311ca2a,open_n69}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b8581517 (
    .a(al_11033702[48]),
    .b(1'b0),
    .c(al_1311ca2a),
    .o({al_cc41fd76,open_n70}));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_affc23c8 (
    .a(numerator[0]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[0]),
    .e(al_c67bebad[0]),
    .o(al_9bfb1470[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_7e4247d5 (
    .a(numerator[10]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[10]),
    .e(al_c67bebad[10]),
    .o(al_9bfb1470[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8f76e334 (
    .a(numerator[11]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[11]),
    .e(al_c67bebad[11]),
    .o(al_9bfb1470[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_43c29c9e (
    .a(numerator[12]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[12]),
    .e(al_c67bebad[12]),
    .o(al_9bfb1470[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_dcb75b0 (
    .a(numerator[13]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[13]),
    .e(al_c67bebad[13]),
    .o(al_9bfb1470[13]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_e1773c9b (
    .a(numerator[14]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[14]),
    .e(al_c67bebad[14]),
    .o(al_9bfb1470[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8e3693cb (
    .a(numerator[15]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[15]),
    .e(al_c67bebad[15]),
    .o(al_9bfb1470[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_79948be9 (
    .a(numerator[16]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[16]),
    .e(al_c67bebad[16]),
    .o(al_9bfb1470[16]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_cd0015f2 (
    .a(numerator[17]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[17]),
    .e(al_c67bebad[17]),
    .o(al_9bfb1470[17]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_5eba52cf (
    .a(numerator[18]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[18]),
    .e(al_c67bebad[18]),
    .o(al_9bfb1470[18]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_fd435063 (
    .a(numerator[19]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[19]),
    .e(al_c67bebad[19]),
    .o(al_9bfb1470[19]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_db832082 (
    .a(numerator[1]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[1]),
    .e(al_c67bebad[1]),
    .o(al_9bfb1470[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_e01dd5be (
    .a(numerator[20]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[20]),
    .e(al_c67bebad[20]),
    .o(al_9bfb1470[20]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3caca9c9 (
    .a(numerator[21]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[21]),
    .e(al_c67bebad[21]),
    .o(al_9bfb1470[21]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_daadae89 (
    .a(numerator[22]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[22]),
    .e(al_c67bebad[22]),
    .o(al_9bfb1470[22]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_29e14add (
    .a(numerator[23]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[23]),
    .e(al_c67bebad[23]),
    .o(al_9bfb1470[23]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_144036ec (
    .a(numerator[24]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[24]),
    .e(al_c67bebad[24]),
    .o(al_9bfb1470[24]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b86a6dbf (
    .a(numerator[25]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[25]),
    .e(al_c67bebad[25]),
    .o(al_9bfb1470[25]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_47ac1c09 (
    .a(numerator[26]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[26]),
    .e(al_c67bebad[26]),
    .o(al_9bfb1470[26]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_248ff2e3 (
    .a(numerator[27]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[27]),
    .e(al_c67bebad[27]),
    .o(al_9bfb1470[27]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_f01911bd (
    .a(numerator[28]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[28]),
    .e(al_c67bebad[28]),
    .o(al_9bfb1470[28]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_67954d07 (
    .a(numerator[29]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[29]),
    .e(al_c67bebad[29]),
    .o(al_9bfb1470[29]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3e04c0e7 (
    .a(numerator[2]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[2]),
    .e(al_c67bebad[2]),
    .o(al_9bfb1470[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3cf932bd (
    .a(numerator[30]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[30]),
    .e(al_c67bebad[30]),
    .o(al_9bfb1470[30]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_4e4f5c0d (
    .a(numerator[31]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[31]),
    .e(al_c67bebad[31]),
    .o(al_9bfb1470[31]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b86e3fac (
    .a(numerator[3]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[3]),
    .e(al_c67bebad[3]),
    .o(al_9bfb1470[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_1f499def (
    .a(numerator[4]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[4]),
    .e(al_c67bebad[4]),
    .o(al_9bfb1470[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8f1711f3 (
    .a(numerator[5]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[5]),
    .e(al_c67bebad[5]),
    .o(al_9bfb1470[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_6e1c653d (
    .a(numerator[6]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[6]),
    .e(al_c67bebad[6]),
    .o(al_9bfb1470[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b46e3fd7 (
    .a(numerator[7]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[7]),
    .e(al_c67bebad[7]),
    .o(al_9bfb1470[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d21f8608 (
    .a(numerator[8]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[8]),
    .e(al_c67bebad[8]),
    .o(al_9bfb1470[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_42e41119 (
    .a(numerator[9]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[9]),
    .e(al_c67bebad[9]),
    .o(al_9bfb1470[9]));
  AL_DFF_0 al_b26d62bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_0 al_809f7104 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_0 al_c1468025 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_0 al_c19d8344 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[3]));
  AL_DFF_0 al_ca1eda73 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[4]));
  AL_DFF_0 al_fa89b429 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[5]));
  AL_DFF_0 al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[8]));
  AL_DFF_0 al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[9]));
  AL_DFF_0 al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[10]));
  AL_DFF_0 al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[11]));
  AL_DFF_0 al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[12]));
  AL_DFF_0 al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[13]));
  AL_DFF_0 al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[14]));
  AL_DFF_0 al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[15]));
  AL_DFF_0 al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[16]));
  AL_DFF_0 al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[17]));
  AL_DFF_0 al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[0]));
  AL_DFF_0 al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[18]));
  AL_DFF_0 al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[19]));
  AL_DFF_0 al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[20]));
  AL_DFF_0 al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[21]));
  AL_DFF_0 al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[22]));
  AL_DFF_0 al_5e95843a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[23]));
  AL_DFF_0 al_d701a9b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[24]));
  AL_DFF_0 al_420d26fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[25]));
  AL_DFF_0 al_eb274ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[27]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[26]));
  AL_DFF_0 al_59566ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[28]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[27]));
  AL_DFF_0 al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[1]));
  AL_DFF_0 al_88ac72e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[29]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[28]));
  AL_DFF_0 al_415d213a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[30]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[29]));
  AL_DFF_0 al_2589b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[31]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[30]));
  AL_DFF_0 al_d3625316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[31]));
  AL_DFF_0 al_a773e9fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[32]));
  AL_DFF_0 al_b5a98930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[33]));
  AL_DFF_0 al_84e187a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[34]));
  AL_DFF_0 al_f3095820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[35]));
  AL_DFF_0 al_9b82a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[36]));
  AL_DFF_0 al_e2ab1094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[37]));
  AL_DFF_0 al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[2]));
  AL_DFF_0 al_a247c67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[38]));
  AL_DFF_0 al_538bab61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[39]));
  AL_DFF_0 al_39eff7a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[40]));
  AL_DFF_0 al_da740eac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[41]));
  AL_DFF_0 al_a1f5e6e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[42]));
  AL_DFF_0 al_73905df6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[43]));
  AL_DFF_0 al_7587b9d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[44]));
  AL_DFF_0 al_cb0b2132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[45]));
  AL_DFF_0 al_79136648 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[46]));
  AL_DFF_0 al_a8eb1e63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[47]));
  AL_DFF_0 al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[3]));
  AL_DFF_0 al_b20ad0fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[48]));
  AL_DFF_0 al_6b481302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[49]));
  AL_DFF_0 al_aa48a4a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[50]));
  AL_DFF_0 al_16453eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[51]));
  AL_DFF_0 al_78700b2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[52]));
  AL_DFF_0 al_3ec4517b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[53]));
  AL_DFF_0 al_f742b91d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[54]));
  AL_DFF_0 al_63888a93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[55]));
  AL_DFF_0 al_3da78364 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[56]));
  AL_DFF_0 al_3d3489ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[57]));
  AL_DFF_0 al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[4]));
  AL_DFF_0 al_d5896133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[58]));
  AL_DFF_0 al_6713d36c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[59]));
  AL_DFF_0 al_498618ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[60]));
  AL_DFF_0 al_f25bea6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[61]));
  AL_DFF_0 al_2e792170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[31]),
    .en(1'b1),
    .sr(~start),
    .ss(1'b0),
    .q(al_11033702[62]));
  AL_DFF_0 al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[5]));
  AL_DFF_0 al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[6]));
  AL_DFF_0 al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[7]));
  AL_DFF_0 al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[8]));
  AL_DFF_0 al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[9]));
  AL_DFF_0 al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[10]));
  AL_DFF_0 al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[11]));
  AL_DFF_0 al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[12]));
  AL_DFF_0 al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[13]));
  AL_DFF_0 al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[14]));
  AL_DFF_0 al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[15]));
  AL_DFF_0 al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[16]));
  AL_DFF_0 al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[17]));
  AL_DFF_0 al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[0]));
  AL_DFF_0 al_2149b062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[18]));
  AL_DFF_0 al_56d82898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[19]));
  AL_DFF_0 al_c8bec57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[20]));
  AL_DFF_0 al_1f071837 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[21]));
  AL_DFF_0 al_9acbb644 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[22]));
  AL_DFF_0 al_286bd0de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[23]));
  AL_DFF_0 al_7e8bb9f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[24]));
  AL_DFF_0 al_d4e324dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[25]));
  AL_DFF_0 al_bcaf406d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[26]));
  AL_DFF_0 al_20d194ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[27]));
  AL_DFF_0 al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[1]));
  AL_DFF_0 al_6402198 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[28]));
  AL_DFF_0 al_3f7239b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[29]));
  AL_DFF_0 al_33cd891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[30]));
  AL_DFF_0 al_28b9e853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[31]));
  AL_DFF_0 al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[2]));
  AL_DFF_0 al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[3]));
  AL_DFF_0 al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[4]));
  AL_DFF_0 al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[5]));
  AL_DFF_0 al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[6]));
  AL_DFF_0 al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[7]));
  AL_DFF_0 al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_0 al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_0 al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_0 al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_0 al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_0 al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_0 al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_0 al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_0 al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_0 al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_0 al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_0 al_68082bd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_0 al_d9e8ef9f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_0 al_39169fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_0 al_c179532 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[21]));
  AL_DFF_0 al_7d105784 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[22]));
  AL_DFF_0 al_573a0a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[23]));
  AL_DFF_0 al_d0deffcb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[24]));
  AL_DFF_0 al_150254f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[25]));
  AL_DFF_0 al_47f1ba67 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[26]));
  AL_DFF_0 al_3f6c28d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[27]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[27]));
  AL_DFF_0 al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_0 al_930b6560 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[28]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[28]));
  AL_DFF_0 al_46a886ac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[29]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[29]));
  AL_DFF_0 al_5c18d1b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[30]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[30]));
  AL_DFF_0 al_f94ac09a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[31]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[31]));
  AL_DFF_0 al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_0 al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_0 al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_0 al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_0 al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_0 al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_0 al_ce6e5997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[8]));
  AL_DFF_0 al_7c322425 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[9]));
  AL_DFF_0 al_1f65ec13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[10]));
  AL_DFF_0 al_63457b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[11]));
  AL_DFF_0 al_11fe6cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[12]));
  AL_DFF_0 al_9cfb6f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[13]));
  AL_DFF_0 al_40b705d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[14]));
  AL_DFF_0 al_cbb21b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[15]));
  AL_DFF_0 al_a743530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[16]));
  AL_DFF_0 al_50032887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[17]));
  AL_DFF_0 al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c61b4192),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[0]));
  AL_DFF_0 al_db3b2b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[18]));
  AL_DFF_0 al_4496adb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[19]));
  AL_DFF_0 al_db38e2c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[20]));
  AL_DFF_0 al_b910420c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[21]));
  AL_DFF_0 al_90d7e42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[22]));
  AL_DFF_0 al_f16a60a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[23]));
  AL_DFF_0 al_91adf23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[24]));
  AL_DFF_0 al_77ecd5d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[25]));
  AL_DFF_0 al_149f3658 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[26]));
  AL_DFF_0 al_8734a4b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[27]));
  AL_DFF_0 al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[1]));
  AL_DFF_0 al_5bba43cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[27]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[28]));
  AL_DFF_0 al_505e168f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[28]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[29]));
  AL_DFF_0 al_a288ce99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[29]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[30]));
  AL_DFF_0 al_930333c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[30]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[31]));
  AL_DFF_0 al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[2]));
  AL_DFF_0 al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[3]));
  AL_DFF_0 al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[4]));
  AL_DFF_0 al_e7cc423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[5]));
  AL_DFF_0 al_2c6ea385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[6]));
  AL_DFF_0 al_a356779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[7]));
  AL_DFF_0 al_f27b108d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_0 al_d1a67c2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_0 al_a7f95d18 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_0 al_da9c9cea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_0 al_40fd9462 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[12]));
  AL_DFF_0 al_ac95b5a9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[13]));
  AL_DFF_0 al_1a9bbf3f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[14]));
  AL_DFF_0 al_66512653 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[15]));
  AL_DFF_0 al_ec92959e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[16]));
  AL_DFF_0 al_efe05263 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[17]));
  AL_DFF_0 al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_0 al_79481707 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[18]));
  AL_DFF_0 al_ed94bd54 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[19]));
  AL_DFF_0 al_a15c98bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[20]));
  AL_DFF_0 al_131a28da (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[21]));
  AL_DFF_0 al_73557a1d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[22]));
  AL_DFF_0 al_a7de7e20 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[23]));
  AL_DFF_0 al_4c32dd42 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[24]));
  AL_DFF_0 al_e05106af (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[25]));
  AL_DFF_0 al_2d9f3ce8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[26]));
  AL_DFF_0 al_de36f4d0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[27]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[27]));
  AL_DFF_0 al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_0 al_f763c3ab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[28]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[28]));
  AL_DFF_0 al_f3dc4f4c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[29]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[29]));
  AL_DFF_0 al_d8cfba43 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[30]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[30]));
  AL_DFF_0 al_d6316b06 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[31]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[31]));
  AL_DFF_0 al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_0 al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_0 al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_0 al_2ccbdc6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_0 al_2c62c395 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_0 al_ee1990ef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_1315ed94[7]),
    .b(al_11033702[7]),
    .c(al_7b07bb65),
    .o({al_9df2af8f,al_c67bebad[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_1315ed94[8]),
    .b(al_11033702[8]),
    .c(al_9df2af8f),
    .o({al_df20ca5b,al_c67bebad[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_1315ed94[9]),
    .b(al_11033702[9]),
    .c(al_df20ca5b),
    .o({al_ab6a0e7,al_c67bebad[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_1315ed94[10]),
    .b(al_11033702[10]),
    .c(al_ab6a0e7),
    .o({al_3f047599,al_c67bebad[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_1315ed94[11]),
    .b(al_11033702[11]),
    .c(al_3f047599),
    .o({al_b4d1b2a2,al_c67bebad[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_1315ed94[12]),
    .b(al_11033702[12]),
    .c(al_b4d1b2a2),
    .o({al_469cb985,al_c67bebad[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_1315ed94[13]),
    .b(al_11033702[13]),
    .c(al_469cb985),
    .o({al_ffb568cb,al_c67bebad[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_1315ed94[14]),
    .b(al_11033702[14]),
    .c(al_ffb568cb),
    .o({al_8f0bd67f,al_c67bebad[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_1315ed94[15]),
    .b(al_11033702[15]),
    .c(al_8f0bd67f),
    .o({al_ee5c4865,al_c67bebad[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_1315ed94[16]),
    .b(al_11033702[16]),
    .c(al_ee5c4865),
    .o({al_c617ea0a,al_c67bebad[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_d21ff3d4,open_n73}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_1315ed94[17]),
    .b(al_11033702[17]),
    .c(al_c617ea0a),
    .o({al_c36dd466,al_c67bebad[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_1315ed94[18]),
    .b(al_11033702[18]),
    .c(al_c36dd466),
    .o({al_cbd8eebc,al_c67bebad[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_1315ed94[19]),
    .b(al_11033702[19]),
    .c(al_cbd8eebc),
    .o({al_c8debd9c,al_c67bebad[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_1315ed94[20]),
    .b(al_11033702[20]),
    .c(al_c8debd9c),
    .o({al_73a2ed86,al_c67bebad[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_1315ed94[21]),
    .b(al_11033702[21]),
    .c(al_73a2ed86),
    .o({al_c8a237ee,al_c67bebad[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e359bb16 (
    .a(al_1315ed94[22]),
    .b(al_11033702[22]),
    .c(al_c8a237ee),
    .o({al_2945efc4,al_c67bebad[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6af83b3 (
    .a(al_1315ed94[23]),
    .b(al_11033702[23]),
    .c(al_2945efc4),
    .o({al_a649c440,al_c67bebad[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_717da7cc (
    .a(al_1315ed94[24]),
    .b(al_11033702[24]),
    .c(al_a649c440),
    .o({al_90e69cc8,al_c67bebad[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_916a9569 (
    .a(al_1315ed94[25]),
    .b(al_11033702[25]),
    .c(al_90e69cc8),
    .o({al_25b33d0e,al_c67bebad[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b53f57fa (
    .a(al_1315ed94[26]),
    .b(al_11033702[26]),
    .c(al_25b33d0e),
    .o({al_ea1005e8,al_c67bebad[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_1315ed94[0]),
    .b(al_11033702[0]),
    .c(al_d21ff3d4),
    .o({al_20da7cd1,al_c67bebad[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_edf2dc1f (
    .a(al_1315ed94[27]),
    .b(al_11033702[27]),
    .c(al_ea1005e8),
    .o({al_128ecb61,al_c67bebad[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a98a3ed7 (
    .a(al_1315ed94[28]),
    .b(al_11033702[28]),
    .c(al_128ecb61),
    .o({al_fb8ac41d,al_c67bebad[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_168d24d3 (
    .a(al_1315ed94[29]),
    .b(al_11033702[29]),
    .c(al_fb8ac41d),
    .o({al_f6cfbe3c,al_c67bebad[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c524c75b (
    .a(al_1315ed94[30]),
    .b(al_11033702[30]),
    .c(al_f6cfbe3c),
    .o({al_ec2ed332,al_c67bebad[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86f90ba9 (
    .a(al_1315ed94[31]),
    .b(al_11033702[31]),
    .c(al_ec2ed332),
    .o({open_n74,al_c67bebad[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_1315ed94[1]),
    .b(al_11033702[1]),
    .c(al_20da7cd1),
    .o({al_4b6c2990,al_c67bebad[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_1315ed94[2]),
    .b(al_11033702[2]),
    .c(al_4b6c2990),
    .o({al_2a9315a6,al_c67bebad[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_1315ed94[3]),
    .b(al_11033702[3]),
    .c(al_2a9315a6),
    .o({al_b9c5d958,al_c67bebad[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_1315ed94[4]),
    .b(al_11033702[4]),
    .c(al_b9c5d958),
    .o({al_56630a35,al_c67bebad[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_1315ed94[5]),
    .b(al_11033702[5]),
    .c(al_56630a35),
    .o({al_a1b0b17a,al_c67bebad[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_1315ed94[6]),
    .b(al_11033702[6]),
    .c(al_a1b0b17a),
    .o({al_7b07bb65,al_c67bebad[6]}));

endmodule 

