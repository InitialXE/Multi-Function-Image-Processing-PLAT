// Verilog netlist created by Tang Dynasty v5.6.119222
// Sat Oct 19 17:02:15 2024

`timescale 1ns / 1ps
module Diver_64
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [63:0] denominator;
  input [63:0] numerator;
  input rst;
  input start;
  output done;
  output [63:0] quotient;
  output [63:0] remainder;

  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 64;
  parameter W_NUM = 64;
  // localparam W_CNT = 7;
  wire [6:0] al_1deac949;
  wire [6:0] al_d0dc52fd;
  wire [6:0] al_537e4616;
  wire [126:0] al_11033702;
  wire [126:0] al_1c1b24e7;
  wire [63:0] al_1315ed94;
  wire [63:0] al_9bfb1470;
  wire [126:0] al_c67bebad;
  wire [63:0] al_327525b3;
  wire al_a707256f;
  wire al_92580e69;
  wire al_ee343458;
  wire al_556ce633;
  wire al_aefd8b68;
  wire al_32ed25d3;
  wire al_2fcc6939;
  wire al_9673d977;
  wire al_a9fbe072;
  wire al_3973d008;
  wire al_4c40b6e5;
  wire al_d63e42fe;
  wire al_b4fc1000;
  wire al_ab829401;
  wire al_b7ca2ed;
  wire al_22a7ce9f;
  wire al_f5902502;
  wire al_b83a67b2;
  wire al_540b209;
  wire al_27e1f3bc;
  wire al_e64e5f1c;
  wire al_e761a920;
  wire al_42ead886;
  wire al_f5a327ab;
  wire al_b23e28b5;
  wire al_283f8d98;
  wire al_516747bd;
  wire al_88a2e01;
  wire al_424d2e3a;
  wire al_5d3a435a;
  wire al_4a5ad68f;
  wire al_9646e713;
  wire al_6cee34b4;
  wire al_9015d2c4;
  wire al_64efb4d0;
  wire al_2d9efd6f;
  wire al_e033469;
  wire al_52f68b55;
  wire al_6b2ca00d;
  wire al_92782c7;
  wire al_ba378049;
  wire al_abb07f01;
  wire al_3a3b377;
  wire al_f762b252;
  wire al_6c2df81c;
  wire al_81606498;
  wire al_fef7e453;
  wire al_84e7266e;
  wire al_5866a5aa;
  wire al_18356e63;
  wire al_4bbb767a;
  wire al_5b37f318;
  wire al_19d272d0;
  wire al_7a6c3f49;
  wire al_59d0e94d;
  wire al_1311ca2a;
  wire al_cc41fd76;
  wire al_9d116ec6;
  wire al_31a76718;
  wire al_728d165d;
  wire al_3c978099;
  wire al_806cd1d1;
  wire al_21e6aa37;
  wire al_d47fc616;
  wire al_a4c56fd2;
  wire al_3aecfb13;
  wire al_a04afdc3;
  wire al_c8596675;
  wire al_26fbd6b;
  wire al_98b263c2;
  wire al_973a6162;
  wire al_7f705d1c;
  wire al_3e979242;
  wire al_73e89f8d;
  wire al_3e495ddf;
  wire al_967c3147;
  wire al_a8cd9f86;
  wire al_79fd50f4;
  wire al_dea4bcb5;
  wire al_ebbda417;
  wire al_36d61c73;
  wire al_fc799980;
  wire al_61806561;
  wire al_d6e4269b;
  wire al_83952368;
  wire al_d433e354;
  wire al_2720c153;
  wire al_b608a891;
  wire al_c18afe64;
  wire al_43e46bab;
  wire al_deee90f;
  wire al_b33d810f;
  wire al_76566ccb;
  wire al_62f0e636;
  wire al_313f5eb8;
  wire al_3d87e86;
  wire al_6fdd3f2c;
  wire al_a7ae70d9;
  wire al_1cb30711;
  wire al_a5d67dd;
  wire al_47366a3a;
  wire al_b4520bce;
  wire al_83fdc521;
  wire al_6a142be1;
  wire al_886f9b5;
  wire al_c9ddd690;
  wire al_95dff75a;
  wire al_4fb90b24;
  wire al_d2bb56b2;
  wire al_18212275;
  wire al_48eda8fd;
  wire al_75eb6ef4;
  wire al_95d30237;
  wire al_8069d0e;
  wire al_596b00a4;
  wire al_502a8237;
  wire al_1b1896c0;
  wire al_4d1a7554;
  wire al_453470b8;
  wire al_ef7500a8;
  wire al_c394171a;
  wire al_83dfff25;
  wire al_3b83b50f;
  wire al_577b588f;
  wire al_ead8205b;
  wire al_815e6466;
  wire al_7813b728;
  wire al_e6d09cdc;
  wire al_a99d77d6;
  wire al_36eba989;
  wire al_477dc4b4;
  wire al_f8ec5b6e;
  wire al_3d132403;
  wire al_dcaa6fc2;
  wire al_c9a7f349;
  wire al_bce8a12e;
  wire al_42574dc6;
  wire al_56f6746e;
  wire al_62cc2266;
  wire al_3be447ce;
  wire al_76e76f5;
  wire al_40413c0d;
  wire al_a2e09ed2;
  wire al_ea253fce;
  wire al_f7bb199b;
  wire al_db6717b5;
  wire al_23548cb7;
  wire al_cb050ae2;
  wire al_9fd06da;
  wire al_b855c346;
  wire al_8f42824f;
  wire al_f2495321;
  wire al_c93cd92e;
  wire al_25204b25;
  wire al_293fb40c;
  wire al_9ea96644;
  wire al_256dce3c;
  wire al_541277c5;
  wire al_111d7f99;
  wire al_caa8d207;
  wire al_fc8fe5d7;
  wire al_c7bb362c;
  wire al_664b4df5;
  wire al_17484234;
  wire al_d77280bf;
  wire al_f0d67edc;
  wire al_c2c0e4c3;
  wire al_f9bb2b5f;
  wire al_72bacdf8;
  wire al_494f78de;
  wire al_63d7a2ad;
  wire al_3de4e7;
  wire al_9a3c1ab7;
  wire al_16b85269;
  wire al_38249694;
  wire al_f6144b57;
  wire al_6da3c5cb;
  wire al_996323c0;
  wire al_edd3bfe4;
  wire al_440c7d0a;
  wire al_4629f076;
  wire al_689ae363;
  wire al_d264df46;
  wire al_29fe8473;
  wire al_a0aced5d;
  wire al_bd3178ec;
  wire al_2a30141f;
  wire al_e391dfd4;
  wire al_c31d4d4f;
  wire al_432a2e5b;
  wire al_59ff8a59;
  wire al_c27564f1;
  wire al_dcd01a2d;
  wire al_9d2f5762;
  wire al_7cb87941;
  wire al_5c338988;
  wire al_9040c841;
  wire al_3f505dba;
  wire al_1d0cd6c7;
  wire al_114eba31;
  wire al_c61b4192;
  wire al_b27e69ab;

  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b22ad72b (
    .a(al_1deac949[3]),
    .b(1'b0),
    .c(al_556ce633),
    .o({al_aefd8b68,al_537e4616[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_37642c3c (
    .a(al_1deac949[4]),
    .b(1'b0),
    .c(al_aefd8b68),
    .o({al_32ed25d3,al_537e4616[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a06a895b (
    .a(al_1deac949[5]),
    .b(1'b0),
    .c(al_32ed25d3),
    .o({al_2fcc6939,al_537e4616[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_877fa7f9 (
    .a(al_1deac949[6]),
    .b(1'b0),
    .c(al_2fcc6939),
    .o({open_n0,al_537e4616[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_a4d828f2 (
    .a(1'b0),
    .o({al_a707256f,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8b186716 (
    .a(al_1deac949[0]),
    .b(1'b1),
    .c(al_a707256f),
    .o({al_92580e69,al_537e4616[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3d917c9c (
    .a(al_1deac949[1]),
    .b(1'b0),
    .c(al_92580e69),
    .o({al_ee343458,al_537e4616[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e7664728 (
    .a(al_1deac949[2]),
    .b(1'b0),
    .c(al_ee343458),
    .o({al_556ce633,al_537e4616[2]}));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_dc50342 (
    .a(al_b27e69ab),
    .b(al_1deac949[0]),
    .c(al_1deac949[6]),
    .o(al_114eba31));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(C*~(A*~(E@D))))"),
    .INIT(32'hdcfcfcdc))
    al_f17cd423 (
    .a(al_b27e69ab),
    .b(start),
    .c(al_537e4616[0]),
    .d(al_1deac949[0]),
    .e(al_1deac949[6]),
    .o(al_d0dc52fd[0]));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(A*~(E@D)))"),
    .INIT(32'h10303010))
    al_147e6a1b (
    .a(al_b27e69ab),
    .b(start),
    .c(al_537e4616[1]),
    .d(al_1deac949[0]),
    .e(al_1deac949[6]),
    .o(al_d0dc52fd[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c8620855 (
    .a(start),
    .b(al_537e4616[2]),
    .o(al_d0dc52fd[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6614de08 (
    .a(start),
    .b(al_537e4616[3]),
    .o(al_d0dc52fd[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6dc5f615 (
    .a(start),
    .b(al_537e4616[4]),
    .o(al_d0dc52fd[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_79196817 (
    .a(start),
    .b(al_537e4616[5]),
    .o(al_d0dc52fd[5]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_5e49efe5 (
    .a(al_1deac949[1]),
    .b(al_1deac949[2]),
    .c(al_1deac949[3]),
    .d(al_1deac949[4]),
    .e(al_1deac949[5]),
    .o(al_b27e69ab));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(A*~(E@D)))"),
    .INIT(32'h10303010))
    al_5e91fab8 (
    .a(al_b27e69ab),
    .b(start),
    .c(al_537e4616[6]),
    .d(al_1deac949[0]),
    .e(al_1deac949[6]),
    .o(al_d0dc52fd[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_255fefd8 (
    .a(denominator[37]),
    .b(start),
    .c(al_11033702[101]),
    .o(al_1c1b24e7[100]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_12c563d8 (
    .a(denominator[38]),
    .b(start),
    .c(al_11033702[102]),
    .o(al_1c1b24e7[101]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_104bdaf9 (
    .a(denominator[39]),
    .b(start),
    .c(al_11033702[103]),
    .o(al_1c1b24e7[102]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c9b92492 (
    .a(denominator[40]),
    .b(start),
    .c(al_11033702[104]),
    .o(al_1c1b24e7[103]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_3aa0ca8 (
    .a(denominator[41]),
    .b(start),
    .c(al_11033702[105]),
    .o(al_1c1b24e7[104]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_35cb8410 (
    .a(denominator[42]),
    .b(start),
    .c(al_11033702[106]),
    .o(al_1c1b24e7[105]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cb87df28 (
    .a(denominator[43]),
    .b(start),
    .c(al_11033702[107]),
    .o(al_1c1b24e7[106]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1a92a8e8 (
    .a(denominator[44]),
    .b(start),
    .c(al_11033702[108]),
    .o(al_1c1b24e7[107]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d6f04a44 (
    .a(denominator[45]),
    .b(start),
    .c(al_11033702[109]),
    .o(al_1c1b24e7[108]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_287bd159 (
    .a(denominator[46]),
    .b(start),
    .c(al_11033702[110]),
    .o(al_1c1b24e7[109]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_6c7772dd (
    .a(denominator[47]),
    .b(start),
    .c(al_11033702[111]),
    .o(al_1c1b24e7[110]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8348ab4b (
    .a(denominator[48]),
    .b(start),
    .c(al_11033702[112]),
    .o(al_1c1b24e7[111]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d03f4b0d (
    .a(denominator[49]),
    .b(start),
    .c(al_11033702[113]),
    .o(al_1c1b24e7[112]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_34120f6f (
    .a(denominator[50]),
    .b(start),
    .c(al_11033702[114]),
    .o(al_1c1b24e7[113]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_81a318d6 (
    .a(denominator[51]),
    .b(start),
    .c(al_11033702[115]),
    .o(al_1c1b24e7[114]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_4d5bca5f (
    .a(denominator[52]),
    .b(start),
    .c(al_11033702[116]),
    .o(al_1c1b24e7[115]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7e1bf57c (
    .a(denominator[53]),
    .b(start),
    .c(al_11033702[117]),
    .o(al_1c1b24e7[116]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_eeefb197 (
    .a(denominator[54]),
    .b(start),
    .c(al_11033702[118]),
    .o(al_1c1b24e7[117]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f8190522 (
    .a(denominator[55]),
    .b(start),
    .c(al_11033702[119]),
    .o(al_1c1b24e7[118]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_7761b502 (
    .a(denominator[56]),
    .b(start),
    .c(al_11033702[120]),
    .o(al_1c1b24e7[119]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b1de5487 (
    .a(denominator[57]),
    .b(start),
    .c(al_11033702[121]),
    .o(al_1c1b24e7[120]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_3c3859eb (
    .a(denominator[58]),
    .b(start),
    .c(al_11033702[122]),
    .o(al_1c1b24e7[121]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_723fd0d4 (
    .a(denominator[59]),
    .b(start),
    .c(al_11033702[123]),
    .o(al_1c1b24e7[122]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_19f92fba (
    .a(denominator[60]),
    .b(start),
    .c(al_11033702[124]),
    .o(al_1c1b24e7[123]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_75538e9c (
    .a(denominator[61]),
    .b(start),
    .c(al_11033702[125]),
    .o(al_1c1b24e7[124]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_89399217 (
    .a(denominator[62]),
    .b(start),
    .c(al_11033702[126]),
    .o(al_1c1b24e7[125]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_cb5602ba (
    .a(denominator[0]),
    .b(start),
    .c(al_11033702[64]),
    .o(al_1c1b24e7[63]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_864b0d81 (
    .a(denominator[1]),
    .b(start),
    .c(al_11033702[65]),
    .o(al_1c1b24e7[64]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a785325 (
    .a(denominator[2]),
    .b(start),
    .c(al_11033702[66]),
    .o(al_1c1b24e7[65]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_3208aa3 (
    .a(denominator[3]),
    .b(start),
    .c(al_11033702[67]),
    .o(al_1c1b24e7[66]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_538719ae (
    .a(denominator[4]),
    .b(start),
    .c(al_11033702[68]),
    .o(al_1c1b24e7[67]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_f420e917 (
    .a(denominator[5]),
    .b(start),
    .c(al_11033702[69]),
    .o(al_1c1b24e7[68]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_97af0053 (
    .a(denominator[6]),
    .b(start),
    .c(al_11033702[70]),
    .o(al_1c1b24e7[69]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_169c3164 (
    .a(denominator[7]),
    .b(start),
    .c(al_11033702[71]),
    .o(al_1c1b24e7[70]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_890551f8 (
    .a(denominator[8]),
    .b(start),
    .c(al_11033702[72]),
    .o(al_1c1b24e7[71]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ba401912 (
    .a(denominator[9]),
    .b(start),
    .c(al_11033702[73]),
    .o(al_1c1b24e7[72]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_39a194b8 (
    .a(denominator[10]),
    .b(start),
    .c(al_11033702[74]),
    .o(al_1c1b24e7[73]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b647e30c (
    .a(denominator[11]),
    .b(start),
    .c(al_11033702[75]),
    .o(al_1c1b24e7[74]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_927d24cb (
    .a(denominator[12]),
    .b(start),
    .c(al_11033702[76]),
    .o(al_1c1b24e7[75]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_2c484ba3 (
    .a(denominator[13]),
    .b(start),
    .c(al_11033702[77]),
    .o(al_1c1b24e7[76]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_556d0a36 (
    .a(denominator[14]),
    .b(start),
    .c(al_11033702[78]),
    .o(al_1c1b24e7[77]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_54553297 (
    .a(denominator[15]),
    .b(start),
    .c(al_11033702[79]),
    .o(al_1c1b24e7[78]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_54ee4e80 (
    .a(denominator[16]),
    .b(start),
    .c(al_11033702[80]),
    .o(al_1c1b24e7[79]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_32497269 (
    .a(denominator[17]),
    .b(start),
    .c(al_11033702[81]),
    .o(al_1c1b24e7[80]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_320b31bd (
    .a(denominator[18]),
    .b(start),
    .c(al_11033702[82]),
    .o(al_1c1b24e7[81]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_6d393ce6 (
    .a(denominator[19]),
    .b(start),
    .c(al_11033702[83]),
    .o(al_1c1b24e7[82]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_757696d8 (
    .a(denominator[20]),
    .b(start),
    .c(al_11033702[84]),
    .o(al_1c1b24e7[83]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e984bf1f (
    .a(denominator[21]),
    .b(start),
    .c(al_11033702[85]),
    .o(al_1c1b24e7[84]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_a4693155 (
    .a(denominator[22]),
    .b(start),
    .c(al_11033702[86]),
    .o(al_1c1b24e7[85]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d351bb13 (
    .a(denominator[23]),
    .b(start),
    .c(al_11033702[87]),
    .o(al_1c1b24e7[86]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_78dbe633 (
    .a(denominator[24]),
    .b(start),
    .c(al_11033702[88]),
    .o(al_1c1b24e7[87]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e0fef712 (
    .a(denominator[25]),
    .b(start),
    .c(al_11033702[89]),
    .o(al_1c1b24e7[88]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_575d9281 (
    .a(denominator[26]),
    .b(start),
    .c(al_11033702[90]),
    .o(al_1c1b24e7[89]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ee65dd15 (
    .a(denominator[27]),
    .b(start),
    .c(al_11033702[91]),
    .o(al_1c1b24e7[90]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e197cd2d (
    .a(denominator[28]),
    .b(start),
    .c(al_11033702[92]),
    .o(al_1c1b24e7[91]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8ae9638d (
    .a(denominator[29]),
    .b(start),
    .c(al_11033702[93]),
    .o(al_1c1b24e7[92]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_57b1111a (
    .a(denominator[30]),
    .b(start),
    .c(al_11033702[94]),
    .o(al_1c1b24e7[93]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_6c476d04 (
    .a(denominator[31]),
    .b(start),
    .c(al_11033702[95]),
    .o(al_1c1b24e7[94]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_76ad634e (
    .a(denominator[32]),
    .b(start),
    .c(al_11033702[96]),
    .o(al_1c1b24e7[95]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_65a8159c (
    .a(denominator[33]),
    .b(start),
    .c(al_11033702[97]),
    .o(al_1c1b24e7[96]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_6a1b2120 (
    .a(denominator[34]),
    .b(start),
    .c(al_11033702[98]),
    .o(al_1c1b24e7[97]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_39c4877b (
    .a(denominator[35]),
    .b(start),
    .c(al_11033702[99]),
    .o(al_1c1b24e7[98]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8942d328 (
    .a(denominator[36]),
    .b(start),
    .c(al_11033702[100]),
    .o(al_1c1b24e7[99]));
  AL_DFF_0 al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_114eba31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    al_2c0796e5 (
    .a(1'b1),
    .o({al_9673d977,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c203f32c (
    .a(al_11033702[4]),
    .b(al_1315ed94[4]),
    .c(al_d63e42fe),
    .o({al_b4fc1000,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_32e253fa (
    .a(al_11033702[49]),
    .b(al_1315ed94[49]),
    .c(al_cc41fd76),
    .o({al_9d116ec6,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_17283bfe (
    .a(al_11033702[50]),
    .b(al_1315ed94[50]),
    .c(al_9d116ec6),
    .o({al_31a76718,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_99897af (
    .a(al_11033702[51]),
    .b(al_1315ed94[51]),
    .c(al_31a76718),
    .o({al_728d165d,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_393be1f9 (
    .a(al_11033702[52]),
    .b(al_1315ed94[52]),
    .c(al_728d165d),
    .o({al_3c978099,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_51bcba86 (
    .a(al_11033702[53]),
    .b(al_1315ed94[53]),
    .c(al_3c978099),
    .o({al_806cd1d1,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4193e874 (
    .a(al_11033702[54]),
    .b(al_1315ed94[54]),
    .c(al_806cd1d1),
    .o({al_21e6aa37,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3eaf5f9c (
    .a(al_11033702[55]),
    .b(al_1315ed94[55]),
    .c(al_21e6aa37),
    .o({al_d47fc616,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c5566d1d (
    .a(al_11033702[56]),
    .b(al_1315ed94[56]),
    .c(al_d47fc616),
    .o({al_a4c56fd2,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9eddbd1b (
    .a(al_11033702[57]),
    .b(al_1315ed94[57]),
    .c(al_a4c56fd2),
    .o({al_3aecfb13,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_245f999 (
    .a(al_11033702[58]),
    .b(al_1315ed94[58]),
    .c(al_3aecfb13),
    .o({al_a04afdc3,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_5a2e66a8 (
    .a(al_11033702[5]),
    .b(al_1315ed94[5]),
    .c(al_b4fc1000),
    .o({al_ab829401,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e21d4825 (
    .a(al_11033702[59]),
    .b(al_1315ed94[59]),
    .c(al_a04afdc3),
    .o({al_c8596675,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ef5c91b6 (
    .a(al_11033702[60]),
    .b(al_1315ed94[60]),
    .c(al_c8596675),
    .o({al_26fbd6b,open_n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b2778311 (
    .a(al_11033702[61]),
    .b(al_1315ed94[61]),
    .c(al_26fbd6b),
    .o({al_98b263c2,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ae943c46 (
    .a(al_11033702[62]),
    .b(al_1315ed94[62]),
    .c(al_98b263c2),
    .o({al_973a6162,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_303727b2 (
    .a(al_11033702[63]),
    .b(al_1315ed94[63]),
    .c(al_973a6162),
    .o({al_7f705d1c,open_n23}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b4261c8b (
    .a(al_11033702[64]),
    .b(1'b0),
    .c(al_7f705d1c),
    .o({al_3e979242,open_n24}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_d835addd (
    .a(al_11033702[65]),
    .b(1'b0),
    .c(al_3e979242),
    .o({al_73e89f8d,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8e95838c (
    .a(al_11033702[66]),
    .b(1'b0),
    .c(al_73e89f8d),
    .o({al_3e495ddf,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8bd8b026 (
    .a(al_11033702[67]),
    .b(1'b0),
    .c(al_3e495ddf),
    .o({al_967c3147,open_n27}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_5cebd753 (
    .a(al_11033702[68]),
    .b(1'b0),
    .c(al_967c3147),
    .o({al_a8cd9f86,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_2f287d12 (
    .a(al_11033702[6]),
    .b(al_1315ed94[6]),
    .c(al_ab829401),
    .o({al_b7ca2ed,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a5d68dd (
    .a(al_11033702[69]),
    .b(1'b0),
    .c(al_a8cd9f86),
    .o({al_79fd50f4,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_6856957b (
    .a(al_11033702[70]),
    .b(1'b0),
    .c(al_79fd50f4),
    .o({al_dea4bcb5,open_n31}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_467b2830 (
    .a(al_11033702[71]),
    .b(1'b0),
    .c(al_dea4bcb5),
    .o({al_ebbda417,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e20a15a0 (
    .a(al_11033702[72]),
    .b(1'b0),
    .c(al_ebbda417),
    .o({al_36d61c73,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1c6872f7 (
    .a(al_11033702[73]),
    .b(1'b0),
    .c(al_36d61c73),
    .o({al_fc799980,open_n34}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_43fa004d (
    .a(al_11033702[74]),
    .b(1'b0),
    .c(al_fc799980),
    .o({al_61806561,open_n35}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_7c2c34f1 (
    .a(al_11033702[75]),
    .b(1'b0),
    .c(al_61806561),
    .o({al_d6e4269b,open_n36}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_bc1c79b (
    .a(al_11033702[76]),
    .b(1'b0),
    .c(al_d6e4269b),
    .o({al_83952368,open_n37}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8e174ca (
    .a(al_11033702[77]),
    .b(1'b0),
    .c(al_83952368),
    .o({al_d433e354,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_635a03cd (
    .a(al_11033702[78]),
    .b(1'b0),
    .c(al_d433e354),
    .o({al_2720c153,open_n39}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9ce86edd (
    .a(al_11033702[7]),
    .b(al_1315ed94[7]),
    .c(al_b7ca2ed),
    .o({al_22a7ce9f,open_n40}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_2ea0249a (
    .a(al_11033702[79]),
    .b(1'b0),
    .c(al_2720c153),
    .o({al_b608a891,open_n41}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1f2c5492 (
    .a(al_11033702[80]),
    .b(1'b0),
    .c(al_b608a891),
    .o({al_c18afe64,open_n42}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_bee70476 (
    .a(al_11033702[81]),
    .b(1'b0),
    .c(al_c18afe64),
    .o({al_43e46bab,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_7db047cb (
    .a(al_11033702[82]),
    .b(1'b0),
    .c(al_43e46bab),
    .o({al_deee90f,open_n44}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_35b152f8 (
    .a(al_11033702[83]),
    .b(1'b0),
    .c(al_deee90f),
    .o({al_b33d810f,open_n45}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b0d23418 (
    .a(al_11033702[84]),
    .b(1'b0),
    .c(al_b33d810f),
    .o({al_76566ccb,open_n46}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_87e836fc (
    .a(al_11033702[85]),
    .b(1'b0),
    .c(al_76566ccb),
    .o({al_62f0e636,open_n47}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1e2cee47 (
    .a(al_11033702[86]),
    .b(1'b0),
    .c(al_62f0e636),
    .o({al_313f5eb8,open_n48}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_2e6eec3 (
    .a(al_11033702[87]),
    .b(1'b0),
    .c(al_313f5eb8),
    .o({al_3d87e86,open_n49}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_6650abde (
    .a(al_11033702[88]),
    .b(1'b0),
    .c(al_3d87e86),
    .o({al_6fdd3f2c,open_n50}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_29f6525 (
    .a(al_11033702[8]),
    .b(al_1315ed94[8]),
    .c(al_22a7ce9f),
    .o({al_f5902502,open_n51}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_994c2245 (
    .a(al_11033702[89]),
    .b(1'b0),
    .c(al_6fdd3f2c),
    .o({al_a7ae70d9,open_n52}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_7772812b (
    .a(al_11033702[90]),
    .b(1'b0),
    .c(al_a7ae70d9),
    .o({al_1cb30711,open_n53}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1bcd7325 (
    .a(al_11033702[91]),
    .b(1'b0),
    .c(al_1cb30711),
    .o({al_a5d67dd,open_n54}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f345e8a7 (
    .a(al_11033702[92]),
    .b(1'b0),
    .c(al_a5d67dd),
    .o({al_47366a3a,open_n55}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ea25c0d7 (
    .a(al_11033702[93]),
    .b(1'b0),
    .c(al_47366a3a),
    .o({al_b4520bce,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3fffbcf (
    .a(al_11033702[94]),
    .b(1'b0),
    .c(al_b4520bce),
    .o({al_83fdc521,open_n57}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e14c53bb (
    .a(al_11033702[95]),
    .b(1'b0),
    .c(al_83fdc521),
    .o({al_6a142be1,open_n58}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_26133636 (
    .a(al_11033702[96]),
    .b(1'b0),
    .c(al_6a142be1),
    .o({al_886f9b5,open_n59}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c0bde678 (
    .a(al_11033702[97]),
    .b(1'b0),
    .c(al_886f9b5),
    .o({al_c9ddd690,open_n60}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_6b065bfd (
    .a(al_11033702[98]),
    .b(1'b0),
    .c(al_c9ddd690),
    .o({al_95dff75a,open_n61}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f171b4f4 (
    .a(al_11033702[0]),
    .b(al_1315ed94[0]),
    .c(al_9673d977),
    .o({al_a9fbe072,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e9c7012b (
    .a(al_11033702[9]),
    .b(al_1315ed94[9]),
    .c(al_f5902502),
    .o({al_b83a67b2,open_n63}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4070a54f (
    .a(al_11033702[99]),
    .b(1'b0),
    .c(al_95dff75a),
    .o({al_4fb90b24,open_n64}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_25e866cf (
    .a(al_11033702[100]),
    .b(1'b0),
    .c(al_4fb90b24),
    .o({al_d2bb56b2,open_n65}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4b7cdd77 (
    .a(al_11033702[101]),
    .b(1'b0),
    .c(al_d2bb56b2),
    .o({al_18212275,open_n66}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_47fb2508 (
    .a(al_11033702[102]),
    .b(1'b0),
    .c(al_18212275),
    .o({al_48eda8fd,open_n67}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9898e0dc (
    .a(al_11033702[103]),
    .b(1'b0),
    .c(al_48eda8fd),
    .o({al_75eb6ef4,open_n68}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_25ee9e36 (
    .a(al_11033702[104]),
    .b(1'b0),
    .c(al_75eb6ef4),
    .o({al_95d30237,open_n69}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_39b8c92a (
    .a(al_11033702[105]),
    .b(1'b0),
    .c(al_95d30237),
    .o({al_8069d0e,open_n70}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a00407c1 (
    .a(al_11033702[106]),
    .b(1'b0),
    .c(al_8069d0e),
    .o({al_596b00a4,open_n71}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9314ca10 (
    .a(al_11033702[107]),
    .b(1'b0),
    .c(al_596b00a4),
    .o({al_502a8237,open_n72}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_6b0d0b30 (
    .a(al_11033702[108]),
    .b(1'b0),
    .c(al_502a8237),
    .o({al_1b1896c0,open_n73}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4226b3d1 (
    .a(al_11033702[10]),
    .b(al_1315ed94[10]),
    .c(al_b83a67b2),
    .o({al_540b209,open_n74}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a9827fbf (
    .a(al_11033702[109]),
    .b(1'b0),
    .c(al_1b1896c0),
    .o({al_4d1a7554,open_n75}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ad6e4af7 (
    .a(al_11033702[110]),
    .b(1'b0),
    .c(al_4d1a7554),
    .o({al_453470b8,open_n76}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_5a197faa (
    .a(al_11033702[111]),
    .b(1'b0),
    .c(al_453470b8),
    .o({al_ef7500a8,open_n77}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_11b6f964 (
    .a(al_11033702[112]),
    .b(1'b0),
    .c(al_ef7500a8),
    .o({al_c394171a,open_n78}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_d87bd00d (
    .a(al_11033702[113]),
    .b(1'b0),
    .c(al_c394171a),
    .o({al_83dfff25,open_n79}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_79c960f3 (
    .a(al_11033702[114]),
    .b(1'b0),
    .c(al_83dfff25),
    .o({al_3b83b50f,open_n80}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_38bd56aa (
    .a(al_11033702[115]),
    .b(1'b0),
    .c(al_3b83b50f),
    .o({al_577b588f,open_n81}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_afa09803 (
    .a(al_11033702[116]),
    .b(1'b0),
    .c(al_577b588f),
    .o({al_ead8205b,open_n82}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8d27eafd (
    .a(al_11033702[117]),
    .b(1'b0),
    .c(al_ead8205b),
    .o({al_815e6466,open_n83}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ab6f9a7d (
    .a(al_11033702[118]),
    .b(1'b0),
    .c(al_815e6466),
    .o({al_7813b728,open_n84}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3f6fc47e (
    .a(al_11033702[11]),
    .b(al_1315ed94[11]),
    .c(al_540b209),
    .o({al_27e1f3bc,open_n85}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a88b66c2 (
    .a(al_11033702[119]),
    .b(1'b0),
    .c(al_7813b728),
    .o({al_e6d09cdc,open_n86}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_418d755d (
    .a(al_11033702[120]),
    .b(1'b0),
    .c(al_e6d09cdc),
    .o({al_a99d77d6,open_n87}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4a2a81e2 (
    .a(al_11033702[121]),
    .b(1'b0),
    .c(al_a99d77d6),
    .o({al_36eba989,open_n88}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f5326a41 (
    .a(al_11033702[122]),
    .b(1'b0),
    .c(al_36eba989),
    .o({al_477dc4b4,open_n89}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_876895c5 (
    .a(al_11033702[123]),
    .b(1'b0),
    .c(al_477dc4b4),
    .o({al_f8ec5b6e,open_n90}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a54c39e7 (
    .a(al_11033702[124]),
    .b(1'b0),
    .c(al_f8ec5b6e),
    .o({al_3d132403,open_n91}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_6070900d (
    .a(al_11033702[125]),
    .b(1'b0),
    .c(al_3d132403),
    .o({al_dcaa6fc2,open_n92}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_2ed918ef (
    .a(al_11033702[126]),
    .b(1'b0),
    .c(al_dcaa6fc2),
    .o({al_c9a7f349,open_n93}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4b671a1 (
    .a(1'b0),
    .b(1'b1),
    .c(al_c9a7f349),
    .o({open_n94,al_c61b4192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e17073e0 (
    .a(al_11033702[12]),
    .b(al_1315ed94[12]),
    .c(al_27e1f3bc),
    .o({al_e64e5f1c,open_n95}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ba5a9770 (
    .a(al_11033702[13]),
    .b(al_1315ed94[13]),
    .c(al_e64e5f1c),
    .o({al_e761a920,open_n96}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cb976531 (
    .a(al_11033702[14]),
    .b(al_1315ed94[14]),
    .c(al_e761a920),
    .o({al_42ead886,open_n97}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e5cd5640 (
    .a(al_11033702[15]),
    .b(al_1315ed94[15]),
    .c(al_42ead886),
    .o({al_f5a327ab,open_n98}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e4d1cd55 (
    .a(al_11033702[16]),
    .b(al_1315ed94[16]),
    .c(al_f5a327ab),
    .o({al_b23e28b5,open_n99}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_dc7e8c2c (
    .a(al_11033702[17]),
    .b(al_1315ed94[17]),
    .c(al_b23e28b5),
    .o({al_283f8d98,open_n100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9ed345ca (
    .a(al_11033702[18]),
    .b(al_1315ed94[18]),
    .c(al_283f8d98),
    .o({al_516747bd,open_n101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_441ad9b2 (
    .a(al_11033702[1]),
    .b(al_1315ed94[1]),
    .c(al_a9fbe072),
    .o({al_3973d008,open_n102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_36cc28eb (
    .a(al_11033702[19]),
    .b(al_1315ed94[19]),
    .c(al_516747bd),
    .o({al_88a2e01,open_n103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e18ee10 (
    .a(al_11033702[20]),
    .b(al_1315ed94[20]),
    .c(al_88a2e01),
    .o({al_424d2e3a,open_n104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_99bd7325 (
    .a(al_11033702[21]),
    .b(al_1315ed94[21]),
    .c(al_424d2e3a),
    .o({al_5d3a435a,open_n105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8aa83152 (
    .a(al_11033702[22]),
    .b(al_1315ed94[22]),
    .c(al_5d3a435a),
    .o({al_4a5ad68f,open_n106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1c94cea5 (
    .a(al_11033702[23]),
    .b(al_1315ed94[23]),
    .c(al_4a5ad68f),
    .o({al_9646e713,open_n107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_d0c6e291 (
    .a(al_11033702[24]),
    .b(al_1315ed94[24]),
    .c(al_9646e713),
    .o({al_6cee34b4,open_n108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b1db9e6d (
    .a(al_11033702[25]),
    .b(al_1315ed94[25]),
    .c(al_6cee34b4),
    .o({al_9015d2c4,open_n109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ada8a24f (
    .a(al_11033702[26]),
    .b(al_1315ed94[26]),
    .c(al_9015d2c4),
    .o({al_64efb4d0,open_n110}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_20b06db2 (
    .a(al_11033702[27]),
    .b(al_1315ed94[27]),
    .c(al_64efb4d0),
    .o({al_2d9efd6f,open_n111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cbda5de1 (
    .a(al_11033702[28]),
    .b(al_1315ed94[28]),
    .c(al_2d9efd6f),
    .o({al_e033469,open_n112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9395428b (
    .a(al_11033702[2]),
    .b(al_1315ed94[2]),
    .c(al_3973d008),
    .o({al_4c40b6e5,open_n113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_361a841e (
    .a(al_11033702[29]),
    .b(al_1315ed94[29]),
    .c(al_e033469),
    .o({al_52f68b55,open_n114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a4c08c3d (
    .a(al_11033702[30]),
    .b(al_1315ed94[30]),
    .c(al_52f68b55),
    .o({al_6b2ca00d,open_n115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_d1ded6e4 (
    .a(al_11033702[31]),
    .b(al_1315ed94[31]),
    .c(al_6b2ca00d),
    .o({al_92782c7,open_n116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f71d9d01 (
    .a(al_11033702[32]),
    .b(al_1315ed94[32]),
    .c(al_92782c7),
    .o({al_ba378049,open_n117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_89b6e9ba (
    .a(al_11033702[33]),
    .b(al_1315ed94[33]),
    .c(al_ba378049),
    .o({al_abb07f01,open_n118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_884478e8 (
    .a(al_11033702[34]),
    .b(al_1315ed94[34]),
    .c(al_abb07f01),
    .o({al_3a3b377,open_n119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_160a5400 (
    .a(al_11033702[35]),
    .b(al_1315ed94[35]),
    .c(al_3a3b377),
    .o({al_f762b252,open_n120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ed8ca432 (
    .a(al_11033702[36]),
    .b(al_1315ed94[36]),
    .c(al_f762b252),
    .o({al_6c2df81c,open_n121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8875c6ac (
    .a(al_11033702[37]),
    .b(al_1315ed94[37]),
    .c(al_6c2df81c),
    .o({al_81606498,open_n122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3611ae8a (
    .a(al_11033702[38]),
    .b(al_1315ed94[38]),
    .c(al_81606498),
    .o({al_fef7e453,open_n123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f7ac689a (
    .a(al_11033702[3]),
    .b(al_1315ed94[3]),
    .c(al_4c40b6e5),
    .o({al_d63e42fe,open_n124}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_36e3cff7 (
    .a(al_11033702[39]),
    .b(al_1315ed94[39]),
    .c(al_fef7e453),
    .o({al_84e7266e,open_n125}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c0e0a8b9 (
    .a(al_11033702[40]),
    .b(al_1315ed94[40]),
    .c(al_84e7266e),
    .o({al_5866a5aa,open_n126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1c410bbd (
    .a(al_11033702[41]),
    .b(al_1315ed94[41]),
    .c(al_5866a5aa),
    .o({al_18356e63,open_n127}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b713d9a8 (
    .a(al_11033702[42]),
    .b(al_1315ed94[42]),
    .c(al_18356e63),
    .o({al_4bbb767a,open_n128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cf933874 (
    .a(al_11033702[43]),
    .b(al_1315ed94[43]),
    .c(al_4bbb767a),
    .o({al_5b37f318,open_n129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8a1cf929 (
    .a(al_11033702[44]),
    .b(al_1315ed94[44]),
    .c(al_5b37f318),
    .o({al_19d272d0,open_n130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_732efaa (
    .a(al_11033702[45]),
    .b(al_1315ed94[45]),
    .c(al_19d272d0),
    .o({al_7a6c3f49,open_n131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c7d9970 (
    .a(al_11033702[46]),
    .b(al_1315ed94[46]),
    .c(al_7a6c3f49),
    .o({al_59d0e94d,open_n132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_a1a5dabd (
    .a(al_11033702[47]),
    .b(al_1315ed94[47]),
    .c(al_59d0e94d),
    .o({al_1311ca2a,open_n133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_b8581517 (
    .a(al_11033702[48]),
    .b(al_1315ed94[48]),
    .c(al_1311ca2a),
    .o({al_cc41fd76,open_n134}));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_affc23c8 (
    .a(numerator[0]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[0]),
    .e(al_c67bebad[0]),
    .o(al_9bfb1470[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_7e4247d5 (
    .a(numerator[10]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[10]),
    .e(al_c67bebad[10]),
    .o(al_9bfb1470[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8f76e334 (
    .a(numerator[11]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[11]),
    .e(al_c67bebad[11]),
    .o(al_9bfb1470[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_43c29c9e (
    .a(numerator[12]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[12]),
    .e(al_c67bebad[12]),
    .o(al_9bfb1470[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_dcb75b0 (
    .a(numerator[13]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[13]),
    .e(al_c67bebad[13]),
    .o(al_9bfb1470[13]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_e1773c9b (
    .a(numerator[14]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[14]),
    .e(al_c67bebad[14]),
    .o(al_9bfb1470[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8e3693cb (
    .a(numerator[15]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[15]),
    .e(al_c67bebad[15]),
    .o(al_9bfb1470[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_79948be9 (
    .a(numerator[16]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[16]),
    .e(al_c67bebad[16]),
    .o(al_9bfb1470[16]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_cd0015f2 (
    .a(numerator[17]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[17]),
    .e(al_c67bebad[17]),
    .o(al_9bfb1470[17]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_5eba52cf (
    .a(numerator[18]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[18]),
    .e(al_c67bebad[18]),
    .o(al_9bfb1470[18]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_fd435063 (
    .a(numerator[19]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[19]),
    .e(al_c67bebad[19]),
    .o(al_9bfb1470[19]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_db832082 (
    .a(numerator[1]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[1]),
    .e(al_c67bebad[1]),
    .o(al_9bfb1470[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_e01dd5be (
    .a(numerator[20]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[20]),
    .e(al_c67bebad[20]),
    .o(al_9bfb1470[20]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3caca9c9 (
    .a(numerator[21]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[21]),
    .e(al_c67bebad[21]),
    .o(al_9bfb1470[21]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_daadae89 (
    .a(numerator[22]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[22]),
    .e(al_c67bebad[22]),
    .o(al_9bfb1470[22]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_29e14add (
    .a(numerator[23]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[23]),
    .e(al_c67bebad[23]),
    .o(al_9bfb1470[23]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_144036ec (
    .a(numerator[24]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[24]),
    .e(al_c67bebad[24]),
    .o(al_9bfb1470[24]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b86a6dbf (
    .a(numerator[25]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[25]),
    .e(al_c67bebad[25]),
    .o(al_9bfb1470[25]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_47ac1c09 (
    .a(numerator[26]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[26]),
    .e(al_c67bebad[26]),
    .o(al_9bfb1470[26]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_248ff2e3 (
    .a(numerator[27]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[27]),
    .e(al_c67bebad[27]),
    .o(al_9bfb1470[27]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_f01911bd (
    .a(numerator[28]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[28]),
    .e(al_c67bebad[28]),
    .o(al_9bfb1470[28]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_67954d07 (
    .a(numerator[29]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[29]),
    .e(al_c67bebad[29]),
    .o(al_9bfb1470[29]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3e04c0e7 (
    .a(numerator[2]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[2]),
    .e(al_c67bebad[2]),
    .o(al_9bfb1470[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3cf932bd (
    .a(numerator[30]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[30]),
    .e(al_c67bebad[30]),
    .o(al_9bfb1470[30]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_4e4f5c0d (
    .a(numerator[31]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[31]),
    .e(al_c67bebad[31]),
    .o(al_9bfb1470[31]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_2068acfa (
    .a(numerator[32]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[32]),
    .e(al_c67bebad[32]),
    .o(al_9bfb1470[32]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b3ebb6c2 (
    .a(numerator[33]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[33]),
    .e(al_c67bebad[33]),
    .o(al_9bfb1470[33]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_4b9f6ba7 (
    .a(numerator[34]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[34]),
    .e(al_c67bebad[34]),
    .o(al_9bfb1470[34]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_a50e6b1e (
    .a(numerator[35]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[35]),
    .e(al_c67bebad[35]),
    .o(al_9bfb1470[35]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d603efb8 (
    .a(numerator[36]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[36]),
    .e(al_c67bebad[36]),
    .o(al_9bfb1470[36]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_aa4b1285 (
    .a(numerator[37]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[37]),
    .e(al_c67bebad[37]),
    .o(al_9bfb1470[37]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_dc908fed (
    .a(numerator[38]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[38]),
    .e(al_c67bebad[38]),
    .o(al_9bfb1470[38]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_43edc8aa (
    .a(numerator[39]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[39]),
    .e(al_c67bebad[39]),
    .o(al_9bfb1470[39]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b86e3fac (
    .a(numerator[3]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[3]),
    .e(al_c67bebad[3]),
    .o(al_9bfb1470[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_a9e6fc77 (
    .a(numerator[40]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[40]),
    .e(al_c67bebad[40]),
    .o(al_9bfb1470[40]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_80104e86 (
    .a(numerator[41]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[41]),
    .e(al_c67bebad[41]),
    .o(al_9bfb1470[41]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_660f5106 (
    .a(numerator[42]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[42]),
    .e(al_c67bebad[42]),
    .o(al_9bfb1470[42]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_bafb7113 (
    .a(numerator[43]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[43]),
    .e(al_c67bebad[43]),
    .o(al_9bfb1470[43]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8848ae4b (
    .a(numerator[44]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[44]),
    .e(al_c67bebad[44]),
    .o(al_9bfb1470[44]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d9a7be7a (
    .a(numerator[45]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[45]),
    .e(al_c67bebad[45]),
    .o(al_9bfb1470[45]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_28eb5e48 (
    .a(numerator[46]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[46]),
    .e(al_c67bebad[46]),
    .o(al_9bfb1470[46]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_fd1bc03 (
    .a(numerator[47]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[47]),
    .e(al_c67bebad[47]),
    .o(al_9bfb1470[47]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_edd71546 (
    .a(numerator[48]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[48]),
    .e(al_c67bebad[48]),
    .o(al_9bfb1470[48]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_c9fdf1aa (
    .a(numerator[49]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[49]),
    .e(al_c67bebad[49]),
    .o(al_9bfb1470[49]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_1f499def (
    .a(numerator[4]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[4]),
    .e(al_c67bebad[4]),
    .o(al_9bfb1470[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_4bed6f9d (
    .a(numerator[50]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[50]),
    .e(al_c67bebad[50]),
    .o(al_9bfb1470[50]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d3663408 (
    .a(numerator[51]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[51]),
    .e(al_c67bebad[51]),
    .o(al_9bfb1470[51]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_c9ff37d5 (
    .a(numerator[52]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[52]),
    .e(al_c67bebad[52]),
    .o(al_9bfb1470[52]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_bae4403d (
    .a(numerator[53]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[53]),
    .e(al_c67bebad[53]),
    .o(al_9bfb1470[53]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_bb72e585 (
    .a(numerator[54]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[54]),
    .e(al_c67bebad[54]),
    .o(al_9bfb1470[54]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_9c607d2f (
    .a(numerator[55]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[55]),
    .e(al_c67bebad[55]),
    .o(al_9bfb1470[55]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b0d1e16a (
    .a(numerator[56]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[56]),
    .e(al_c67bebad[56]),
    .o(al_9bfb1470[56]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_52fdfab0 (
    .a(numerator[57]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[57]),
    .e(al_c67bebad[57]),
    .o(al_9bfb1470[57]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_96b2184f (
    .a(numerator[58]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[58]),
    .e(al_c67bebad[58]),
    .o(al_9bfb1470[58]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_ec83fefb (
    .a(numerator[59]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[59]),
    .e(al_c67bebad[59]),
    .o(al_9bfb1470[59]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8f1711f3 (
    .a(numerator[5]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[5]),
    .e(al_c67bebad[5]),
    .o(al_9bfb1470[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d4078049 (
    .a(numerator[60]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[60]),
    .e(al_c67bebad[60]),
    .o(al_9bfb1470[60]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d7599f43 (
    .a(numerator[61]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[61]),
    .e(al_c67bebad[61]),
    .o(al_9bfb1470[61]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_fe8f003f (
    .a(numerator[62]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[62]),
    .e(al_c67bebad[62]),
    .o(al_9bfb1470[62]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_4edaf895 (
    .a(numerator[63]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[63]),
    .e(al_c67bebad[63]),
    .o(al_9bfb1470[63]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_6e1c653d (
    .a(numerator[6]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[6]),
    .e(al_c67bebad[6]),
    .o(al_9bfb1470[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b46e3fd7 (
    .a(numerator[7]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[7]),
    .e(al_c67bebad[7]),
    .o(al_9bfb1470[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d21f8608 (
    .a(numerator[8]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[8]),
    .e(al_c67bebad[8]),
    .o(al_9bfb1470[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_42e41119 (
    .a(numerator[9]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[9]),
    .e(al_c67bebad[9]),
    .o(al_9bfb1470[9]));
  AL_DFF_0 al_b26d62bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_0 al_809f7104 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_0 al_c1468025 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_0 al_c19d8344 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[3]));
  AL_DFF_0 al_ca1eda73 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[4]));
  AL_DFF_0 al_fa89b429 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[5]));
  AL_DFF_0 al_3462fe16 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[6]));
  AL_DFF_0 al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[8]));
  AL_DFF_0 al_1d612f9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[98]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[98]));
  AL_DFF_0 al_606f23d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[99]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[99]));
  AL_DFF_0 al_c4f442ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[100]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[100]));
  AL_DFF_0 al_ce7501a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[101]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[101]));
  AL_DFF_0 al_ce875aed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[102]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[102]));
  AL_DFF_0 al_dbb69d66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[103]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[103]));
  AL_DFF_0 al_81f5861 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[104]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[104]));
  AL_DFF_0 al_f1f27903 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[105]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[105]));
  AL_DFF_0 al_8a0d2848 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[106]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[106]));
  AL_DFF_0 al_64d162c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[107]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[107]));
  AL_DFF_0 al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[9]));
  AL_DFF_0 al_7da5002b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[108]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[108]));
  AL_DFF_0 al_78690025 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[109]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[109]));
  AL_DFF_0 al_4f8d9421 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[110]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[110]));
  AL_DFF_0 al_948b8f4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[111]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[111]));
  AL_DFF_0 al_83aa1770 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[112]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[112]));
  AL_DFF_0 al_ac2f6d59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[113]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[113]));
  AL_DFF_0 al_7c4e2237 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[114]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[114]));
  AL_DFF_0 al_2613b88c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[115]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[115]));
  AL_DFF_0 al_ceda802d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[116]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[116]));
  AL_DFF_0 al_2d135f8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[117]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[117]));
  AL_DFF_0 al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[10]));
  AL_DFF_0 al_61c3fb9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[118]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[118]));
  AL_DFF_0 al_f226845c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[119]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[119]));
  AL_DFF_0 al_586fa12d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[120]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[120]));
  AL_DFF_0 al_f2bad4f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[121]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[121]));
  AL_DFF_0 al_eecaea83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[122]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[122]));
  AL_DFF_0 al_34ccfd1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[123]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[123]));
  AL_DFF_0 al_9ade58dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[124]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[124]));
  AL_DFF_0 al_23580333 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[125]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[125]));
  AL_DFF_0 al_90297b7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[63]),
    .en(1'b1),
    .sr(~start),
    .ss(1'b0),
    .q(al_11033702[126]));
  AL_DFF_0 al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[11]));
  AL_DFF_0 al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[12]));
  AL_DFF_0 al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[13]));
  AL_DFF_0 al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[14]));
  AL_DFF_0 al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[15]));
  AL_DFF_0 al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[16]));
  AL_DFF_0 al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[17]));
  AL_DFF_0 al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[0]));
  AL_DFF_0 al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[18]));
  AL_DFF_0 al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[19]));
  AL_DFF_0 al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[20]));
  AL_DFF_0 al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[21]));
  AL_DFF_0 al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[22]));
  AL_DFF_0 al_5e95843a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[23]));
  AL_DFF_0 al_d701a9b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[24]));
  AL_DFF_0 al_420d26fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[25]));
  AL_DFF_0 al_eb274ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[27]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[26]));
  AL_DFF_0 al_59566ddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[28]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[27]));
  AL_DFF_0 al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[1]));
  AL_DFF_0 al_88ac72e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[29]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[28]));
  AL_DFF_0 al_415d213a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[30]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[29]));
  AL_DFF_0 al_2589b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[31]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[30]));
  AL_DFF_0 al_d3625316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[32]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[31]));
  AL_DFF_0 al_a773e9fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[33]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[32]));
  AL_DFF_0 al_b5a98930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[34]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[33]));
  AL_DFF_0 al_84e187a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[35]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[34]));
  AL_DFF_0 al_f3095820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[36]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[35]));
  AL_DFF_0 al_9b82a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[37]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[36]));
  AL_DFF_0 al_e2ab1094 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[38]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[37]));
  AL_DFF_0 al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[2]));
  AL_DFF_0 al_a247c67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[39]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[38]));
  AL_DFF_0 al_538bab61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[40]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[39]));
  AL_DFF_0 al_39eff7a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[41]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[40]));
  AL_DFF_0 al_da740eac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[42]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[41]));
  AL_DFF_0 al_a1f5e6e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[43]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[42]));
  AL_DFF_0 al_73905df6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[44]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[43]));
  AL_DFF_0 al_7587b9d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[45]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[44]));
  AL_DFF_0 al_cb0b2132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[46]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[45]));
  AL_DFF_0 al_79136648 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[47]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[46]));
  AL_DFF_0 al_a8eb1e63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[48]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[47]));
  AL_DFF_0 al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[3]));
  AL_DFF_0 al_b20ad0fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[49]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[48]));
  AL_DFF_0 al_6b481302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[50]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[49]));
  AL_DFF_0 al_aa48a4a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[51]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[50]));
  AL_DFF_0 al_16453eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[52]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[51]));
  AL_DFF_0 al_78700b2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[53]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[52]));
  AL_DFF_0 al_3ec4517b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[54]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[53]));
  AL_DFF_0 al_f742b91d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[55]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[54]));
  AL_DFF_0 al_63888a93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[56]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[55]));
  AL_DFF_0 al_3da78364 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[57]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[56]));
  AL_DFF_0 al_3d3489ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[58]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[57]));
  AL_DFF_0 al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[4]));
  AL_DFF_0 al_d5896133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[59]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[58]));
  AL_DFF_0 al_6713d36c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[60]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[59]));
  AL_DFF_0 al_498618ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[61]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[60]));
  AL_DFF_0 al_f25bea6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[62]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[61]));
  AL_DFF_0 al_2e792170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[63]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[62]));
  AL_DFF_0 al_10e927f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[63]));
  AL_DFF_0 al_6cdaad66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[64]));
  AL_DFF_0 al_428372bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[65]));
  AL_DFF_0 al_f8209620 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[66]));
  AL_DFF_0 al_96ae94d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[67]));
  AL_DFF_0 al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[5]));
  AL_DFF_0 al_be0c1a24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[68]));
  AL_DFF_0 al_a5d841b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[69]));
  AL_DFF_0 al_b6808dcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[70]));
  AL_DFF_0 al_5fd20133 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[71]));
  AL_DFF_0 al_57550c35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[72]));
  AL_DFF_0 al_a08195e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[73]));
  AL_DFF_0 al_8c7f06d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[74]));
  AL_DFF_0 al_9fa13836 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[75]));
  AL_DFF_0 al_815541d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[76]));
  AL_DFF_0 al_5034b12e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[77]));
  AL_DFF_0 al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[6]));
  AL_DFF_0 al_5620c68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[78]));
  AL_DFF_0 al_45219d16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[79]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[79]));
  AL_DFF_0 al_64a178bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[80]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[80]));
  AL_DFF_0 al_9d8293e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[81]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[81]));
  AL_DFF_0 al_ce49bf1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[82]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[82]));
  AL_DFF_0 al_4fc02135 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[83]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[83]));
  AL_DFF_0 al_3735b737 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[84]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[84]));
  AL_DFF_0 al_e3b5582d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[85]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[85]));
  AL_DFF_0 al_21ceca71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[86]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[86]));
  AL_DFF_0 al_26e3c653 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[87]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[87]));
  AL_DFF_0 al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[7]));
  AL_DFF_0 al_b198e26e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[88]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[88]));
  AL_DFF_0 al_30ff7bbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[89]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[89]));
  AL_DFF_0 al_58f85d1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[90]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[90]));
  AL_DFF_0 al_8c5ed32a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[91]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[91]));
  AL_DFF_0 al_7ac5965 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[92]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[92]));
  AL_DFF_0 al_bd98ac16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[93]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[93]));
  AL_DFF_0 al_cfc49e47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[94]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[94]));
  AL_DFF_0 al_5aef312a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[95]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[95]));
  AL_DFF_0 al_40e1865f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[96]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[96]));
  AL_DFF_0 al_7d0da19f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[97]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[97]));
  AL_DFF_0 al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[8]));
  AL_DFF_0 al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[9]));
  AL_DFF_0 al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[10]));
  AL_DFF_0 al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[11]));
  AL_DFF_0 al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[12]));
  AL_DFF_0 al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[13]));
  AL_DFF_0 al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[14]));
  AL_DFF_0 al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[15]));
  AL_DFF_0 al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[16]));
  AL_DFF_0 al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[17]));
  AL_DFF_0 al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[0]));
  AL_DFF_0 al_2149b062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[18]));
  AL_DFF_0 al_56d82898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[19]));
  AL_DFF_0 al_c8bec57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[20]));
  AL_DFF_0 al_1f071837 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[21]));
  AL_DFF_0 al_9acbb644 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[22]));
  AL_DFF_0 al_286bd0de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[23]));
  AL_DFF_0 al_7e8bb9f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[24]));
  AL_DFF_0 al_d4e324dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[25]));
  AL_DFF_0 al_bcaf406d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[26]));
  AL_DFF_0 al_20d194ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[27]));
  AL_DFF_0 al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[1]));
  AL_DFF_0 al_6402198 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[28]));
  AL_DFF_0 al_3f7239b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[29]));
  AL_DFF_0 al_33cd891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[30]));
  AL_DFF_0 al_28b9e853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[31]));
  AL_DFF_0 al_2da6eeb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[32]));
  AL_DFF_0 al_cca00973 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[33]));
  AL_DFF_0 al_6bc4a040 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[34]));
  AL_DFF_0 al_7cf6bbec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[35]));
  AL_DFF_0 al_3b3f2d26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[36]));
  AL_DFF_0 al_dc5b9d24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[37]));
  AL_DFF_0 al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[2]));
  AL_DFF_0 al_faa19bbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[38]));
  AL_DFF_0 al_33941afe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[39]));
  AL_DFF_0 al_859d7b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[40]));
  AL_DFF_0 al_7f8ef6ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[41]));
  AL_DFF_0 al_efcfba42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[42]));
  AL_DFF_0 al_add7811b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[43]));
  AL_DFF_0 al_f30e50f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[44]));
  AL_DFF_0 al_c8583035 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[45]));
  AL_DFF_0 al_3fc0b4bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[46]));
  AL_DFF_0 al_5d831b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[47]));
  AL_DFF_0 al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[3]));
  AL_DFF_0 al_7b1cfe82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[48]));
  AL_DFF_0 al_41ed5389 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[49]));
  AL_DFF_0 al_a99fa5b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[50]));
  AL_DFF_0 al_84bc2a18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[51]));
  AL_DFF_0 al_f2a3f8de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[52]));
  AL_DFF_0 al_d44591ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[53]));
  AL_DFF_0 al_84f23f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[54]));
  AL_DFF_0 al_c39ae774 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[55]));
  AL_DFF_0 al_5d3fd884 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[56]));
  AL_DFF_0 al_120b5a84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[57]));
  AL_DFF_0 al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[4]));
  AL_DFF_0 al_d54fbc04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[58]));
  AL_DFF_0 al_a1f7f93d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[59]));
  AL_DFF_0 al_b9beab17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[60]));
  AL_DFF_0 al_ac590a10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[61]));
  AL_DFF_0 al_a6976454 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[62]));
  AL_DFF_0 al_c884e8ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[63]));
  AL_DFF_0 al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[5]));
  AL_DFF_0 al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[6]));
  AL_DFF_0 al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[7]));
  AL_DFF_0 al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_0 al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_0 al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_0 al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_0 al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_0 al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_0 al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_0 al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_0 al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_0 al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_0 al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_0 al_68082bd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_0 al_d9e8ef9f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_0 al_39169fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_0 al_c179532 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[21]));
  AL_DFF_0 al_7d105784 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[22]));
  AL_DFF_0 al_573a0a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[23]));
  AL_DFF_0 al_d0deffcb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[24]));
  AL_DFF_0 al_150254f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[25]));
  AL_DFF_0 al_47f1ba67 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[26]));
  AL_DFF_0 al_3f6c28d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[27]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[27]));
  AL_DFF_0 al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_0 al_930b6560 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[28]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[28]));
  AL_DFF_0 al_46a886ac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[29]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[29]));
  AL_DFF_0 al_5c18d1b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[30]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[30]));
  AL_DFF_0 al_f94ac09a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[31]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[31]));
  AL_DFF_0 al_4e65699f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[32]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[32]));
  AL_DFF_0 al_e18c69c7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[33]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[33]));
  AL_DFF_0 al_e1d2b0c2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[34]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[34]));
  AL_DFF_0 al_58830fc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[35]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[35]));
  AL_DFF_0 al_d9d78798 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[36]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[36]));
  AL_DFF_0 al_7013bc9a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[37]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[37]));
  AL_DFF_0 al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_0 al_436ca8bb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[38]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[38]));
  AL_DFF_0 al_4ccfd875 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[39]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[39]));
  AL_DFF_0 al_bb5d438b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[40]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[40]));
  AL_DFF_0 al_3f7dcd40 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[41]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[41]));
  AL_DFF_0 al_c25f43fe (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[42]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[42]));
  AL_DFF_0 al_35c2d44e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[43]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[43]));
  AL_DFF_0 al_f23e3d6c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[44]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[44]));
  AL_DFF_0 al_9df8f24 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[45]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[45]));
  AL_DFF_0 al_d829f573 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[46]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[46]));
  AL_DFF_0 al_2e3b4fdd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[47]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[47]));
  AL_DFF_0 al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_0 al_ec0d726 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[48]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[48]));
  AL_DFF_0 al_97f244c9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[49]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[49]));
  AL_DFF_0 al_567b6740 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[50]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[50]));
  AL_DFF_0 al_31998ccc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[51]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[51]));
  AL_DFF_0 al_a37b1673 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[52]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[52]));
  AL_DFF_0 al_e96a23d8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[53]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[53]));
  AL_DFF_0 al_49894184 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[54]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[54]));
  AL_DFF_0 al_4d71573c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[55]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[55]));
  AL_DFF_0 al_c9a1fd27 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[56]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[56]));
  AL_DFF_0 al_353edd92 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[57]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[57]));
  AL_DFF_0 al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_0 al_33896c84 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[58]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[58]));
  AL_DFF_0 al_372db785 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[59]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[59]));
  AL_DFF_0 al_572f0a39 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[60]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[60]));
  AL_DFF_0 al_6fae33b3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[61]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[61]));
  AL_DFF_0 al_7dabf020 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[62]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[62]));
  AL_DFF_0 al_710039e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[63]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[63]));
  AL_DFF_0 al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_0 al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_0 al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_0 al_ce6e5997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[8]));
  AL_DFF_0 al_7c322425 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[9]));
  AL_DFF_0 al_1f65ec13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[10]));
  AL_DFF_0 al_63457b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[11]));
  AL_DFF_0 al_11fe6cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[12]));
  AL_DFF_0 al_9cfb6f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[13]));
  AL_DFF_0 al_40b705d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[14]));
  AL_DFF_0 al_cbb21b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[15]));
  AL_DFF_0 al_a743530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[16]));
  AL_DFF_0 al_50032887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[17]));
  AL_DFF_0 al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c61b4192),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[0]));
  AL_DFF_0 al_db3b2b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[18]));
  AL_DFF_0 al_4496adb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[18]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[19]));
  AL_DFF_0 al_db38e2c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[19]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[20]));
  AL_DFF_0 al_b910420c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[20]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[21]));
  AL_DFF_0 al_90d7e42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[21]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[22]));
  AL_DFF_0 al_f16a60a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[22]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[23]));
  AL_DFF_0 al_91adf23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[23]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[24]));
  AL_DFF_0 al_77ecd5d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[24]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[25]));
  AL_DFF_0 al_149f3658 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[25]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[26]));
  AL_DFF_0 al_8734a4b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[26]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[27]));
  AL_DFF_0 al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[1]));
  AL_DFF_0 al_5bba43cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[27]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[28]));
  AL_DFF_0 al_505e168f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[28]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[29]));
  AL_DFF_0 al_a288ce99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[29]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[30]));
  AL_DFF_0 al_930333c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[30]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[31]));
  AL_DFF_0 al_5d27e954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[31]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[32]));
  AL_DFF_0 al_f0da03a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[32]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[33]));
  AL_DFF_0 al_c8a0e628 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[33]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[34]));
  AL_DFF_0 al_f689feb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[34]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[35]));
  AL_DFF_0 al_27f9e709 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[35]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[36]));
  AL_DFF_0 al_28d079d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[36]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[37]));
  AL_DFF_0 al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[2]));
  AL_DFF_0 al_be3e1444 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[37]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[38]));
  AL_DFF_0 al_79186d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[38]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[39]));
  AL_DFF_0 al_8a46cd85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[39]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[40]));
  AL_DFF_0 al_aa53ffe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[40]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[41]));
  AL_DFF_0 al_4203609d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[41]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[42]));
  AL_DFF_0 al_40bed0ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[42]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[43]));
  AL_DFF_0 al_ef773c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[43]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[44]));
  AL_DFF_0 al_715ce79a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[44]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[45]));
  AL_DFF_0 al_a733a01f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[45]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[46]));
  AL_DFF_0 al_97115bd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[46]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[47]));
  AL_DFF_0 al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[3]));
  AL_DFF_0 al_da8ba34a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[47]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[48]));
  AL_DFF_0 al_bf47b81b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[48]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[49]));
  AL_DFF_0 al_23770100 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[49]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[50]));
  AL_DFF_0 al_1b3e581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[50]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[51]));
  AL_DFF_0 al_91d20b98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[51]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[52]));
  AL_DFF_0 al_c19fc14a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[52]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[53]));
  AL_DFF_0 al_7e937ee9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[53]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[54]));
  AL_DFF_0 al_78832841 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[54]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[55]));
  AL_DFF_0 al_554bb008 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[55]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[56]));
  AL_DFF_0 al_3726609a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[56]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[57]));
  AL_DFF_0 al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[4]));
  AL_DFF_0 al_6ee699e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[57]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[58]));
  AL_DFF_0 al_e6a6006b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[58]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[59]));
  AL_DFF_0 al_2f20e43d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[59]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[60]));
  AL_DFF_0 al_7e6d452f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[60]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[61]));
  AL_DFF_0 al_36b1076e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[61]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[62]));
  AL_DFF_0 al_3a8f6c9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[62]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[63]));
  AL_DFF_0 al_e7cc423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[5]));
  AL_DFF_0 al_2c6ea385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[6]));
  AL_DFF_0 al_a356779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[7]));
  AL_DFF_0 al_f27b108d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_0 al_d1a67c2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_0 al_a7f95d18 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_0 al_da9c9cea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_0 al_40fd9462 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[12]));
  AL_DFF_0 al_ac95b5a9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[13]));
  AL_DFF_0 al_1a9bbf3f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[14]));
  AL_DFF_0 al_66512653 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[15]));
  AL_DFF_0 al_ec92959e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[16]));
  AL_DFF_0 al_efe05263 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[17]));
  AL_DFF_0 al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_0 al_79481707 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[18]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[18]));
  AL_DFF_0 al_ed94bd54 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[19]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[19]));
  AL_DFF_0 al_a15c98bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[20]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[20]));
  AL_DFF_0 al_131a28da (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[21]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[21]));
  AL_DFF_0 al_73557a1d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[22]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[22]));
  AL_DFF_0 al_a7de7e20 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[23]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[23]));
  AL_DFF_0 al_4c32dd42 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[24]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[24]));
  AL_DFF_0 al_e05106af (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[25]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[25]));
  AL_DFF_0 al_2d9f3ce8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[26]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[26]));
  AL_DFF_0 al_de36f4d0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[27]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[27]));
  AL_DFF_0 al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_0 al_f763c3ab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[28]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[28]));
  AL_DFF_0 al_f3dc4f4c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[29]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[29]));
  AL_DFF_0 al_d8cfba43 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[30]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[30]));
  AL_DFF_0 al_d6316b06 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[31]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[31]));
  AL_DFF_0 al_8cc9cf1e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[32]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[32]));
  AL_DFF_0 al_727888e7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[33]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[33]));
  AL_DFF_0 al_42457074 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[34]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[34]));
  AL_DFF_0 al_a25b8e32 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[35]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[35]));
  AL_DFF_0 al_94674763 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[36]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[36]));
  AL_DFF_0 al_be3f394b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[37]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[37]));
  AL_DFF_0 al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_0 al_4f9b8bbb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[38]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[38]));
  AL_DFF_0 al_c826e53b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[39]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[39]));
  AL_DFF_0 al_88059fd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[40]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[40]));
  AL_DFF_0 al_1923cba2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[41]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[41]));
  AL_DFF_0 al_aa6bee0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[42]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[42]));
  AL_DFF_0 al_ddc7f719 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[43]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[43]));
  AL_DFF_0 al_e224f457 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[44]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[44]));
  AL_DFF_0 al_105930e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[45]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[45]));
  AL_DFF_0 al_4d1b18fa (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[46]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[46]));
  AL_DFF_0 al_8a94269f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[47]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[47]));
  AL_DFF_0 al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_0 al_26e720bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[48]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[48]));
  AL_DFF_0 al_f593af7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[49]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[49]));
  AL_DFF_0 al_9640e362 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[50]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[50]));
  AL_DFF_0 al_4a1cc6f1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[51]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[51]));
  AL_DFF_0 al_2eaa27c5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[52]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[52]));
  AL_DFF_0 al_cc18654a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[53]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[53]));
  AL_DFF_0 al_ff32a167 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[54]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[54]));
  AL_DFF_0 al_ef696938 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[55]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[55]));
  AL_DFF_0 al_348960a3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[56]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[56]));
  AL_DFF_0 al_61e14f5a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[57]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[57]));
  AL_DFF_0 al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_0 al_215cc356 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[58]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[58]));
  AL_DFF_0 al_e8103154 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[59]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[59]));
  AL_DFF_0 al_7ccc43c6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[60]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[60]));
  AL_DFF_0 al_af329b80 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[61]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[61]));
  AL_DFF_0 al_9fff6f0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[62]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[62]));
  AL_DFF_0 al_9f78ce64 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[63]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[63]));
  AL_DFF_0 al_2ccbdc6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_0 al_2c62c395 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_0 al_ee1990ef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_1315ed94[7]),
    .b(al_11033702[7]),
    .c(al_a2e09ed2),
    .o({al_ea253fce,al_c67bebad[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_1315ed94[8]),
    .b(al_11033702[8]),
    .c(al_ea253fce),
    .o({al_f7bb199b,al_c67bebad[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_1315ed94[9]),
    .b(al_11033702[9]),
    .c(al_f7bb199b),
    .o({al_db6717b5,al_c67bebad[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_1315ed94[10]),
    .b(al_11033702[10]),
    .c(al_db6717b5),
    .o({al_23548cb7,al_c67bebad[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_1315ed94[11]),
    .b(al_11033702[11]),
    .c(al_23548cb7),
    .o({al_cb050ae2,al_c67bebad[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_1315ed94[12]),
    .b(al_11033702[12]),
    .c(al_cb050ae2),
    .o({al_9fd06da,al_c67bebad[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_1315ed94[13]),
    .b(al_11033702[13]),
    .c(al_9fd06da),
    .o({al_b855c346,al_c67bebad[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_1315ed94[14]),
    .b(al_11033702[14]),
    .c(al_b855c346),
    .o({al_8f42824f,al_c67bebad[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_1315ed94[15]),
    .b(al_11033702[15]),
    .c(al_8f42824f),
    .o({al_f2495321,al_c67bebad[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_1315ed94[16]),
    .b(al_11033702[16]),
    .c(al_f2495321),
    .o({al_c93cd92e,al_c67bebad[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_bce8a12e,open_n137}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_1315ed94[17]),
    .b(al_11033702[17]),
    .c(al_c93cd92e),
    .o({al_25204b25,al_c67bebad[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_1315ed94[18]),
    .b(al_11033702[18]),
    .c(al_25204b25),
    .o({al_293fb40c,al_c67bebad[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_1315ed94[19]),
    .b(al_11033702[19]),
    .c(al_293fb40c),
    .o({al_9ea96644,al_c67bebad[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_1315ed94[20]),
    .b(al_11033702[20]),
    .c(al_9ea96644),
    .o({al_256dce3c,al_c67bebad[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_1315ed94[21]),
    .b(al_11033702[21]),
    .c(al_256dce3c),
    .o({al_541277c5,al_c67bebad[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e359bb16 (
    .a(al_1315ed94[22]),
    .b(al_11033702[22]),
    .c(al_541277c5),
    .o({al_111d7f99,al_c67bebad[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6af83b3 (
    .a(al_1315ed94[23]),
    .b(al_11033702[23]),
    .c(al_111d7f99),
    .o({al_caa8d207,al_c67bebad[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_717da7cc (
    .a(al_1315ed94[24]),
    .b(al_11033702[24]),
    .c(al_caa8d207),
    .o({al_fc8fe5d7,al_c67bebad[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_916a9569 (
    .a(al_1315ed94[25]),
    .b(al_11033702[25]),
    .c(al_fc8fe5d7),
    .o({al_c7bb362c,al_c67bebad[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b53f57fa (
    .a(al_1315ed94[26]),
    .b(al_11033702[26]),
    .c(al_c7bb362c),
    .o({al_664b4df5,al_c67bebad[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_1315ed94[0]),
    .b(al_11033702[0]),
    .c(al_bce8a12e),
    .o({al_42574dc6,al_c67bebad[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_edf2dc1f (
    .a(al_1315ed94[27]),
    .b(al_11033702[27]),
    .c(al_664b4df5),
    .o({al_17484234,al_c67bebad[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a98a3ed7 (
    .a(al_1315ed94[28]),
    .b(al_11033702[28]),
    .c(al_17484234),
    .o({al_d77280bf,al_c67bebad[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_168d24d3 (
    .a(al_1315ed94[29]),
    .b(al_11033702[29]),
    .c(al_d77280bf),
    .o({al_f0d67edc,al_c67bebad[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c524c75b (
    .a(al_1315ed94[30]),
    .b(al_11033702[30]),
    .c(al_f0d67edc),
    .o({al_c2c0e4c3,al_c67bebad[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86f90ba9 (
    .a(al_1315ed94[31]),
    .b(al_11033702[31]),
    .c(al_c2c0e4c3),
    .o({al_f9bb2b5f,al_c67bebad[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_344fb63e (
    .a(al_1315ed94[32]),
    .b(al_11033702[32]),
    .c(al_f9bb2b5f),
    .o({al_72bacdf8,al_c67bebad[32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fafc8f53 (
    .a(al_1315ed94[33]),
    .b(al_11033702[33]),
    .c(al_72bacdf8),
    .o({al_494f78de,al_c67bebad[33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33de60a (
    .a(al_1315ed94[34]),
    .b(al_11033702[34]),
    .c(al_494f78de),
    .o({al_63d7a2ad,al_c67bebad[34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ae4de70 (
    .a(al_1315ed94[35]),
    .b(al_11033702[35]),
    .c(al_63d7a2ad),
    .o({al_3de4e7,al_c67bebad[35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff46470e (
    .a(al_1315ed94[36]),
    .b(al_11033702[36]),
    .c(al_3de4e7),
    .o({al_9a3c1ab7,al_c67bebad[36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_1315ed94[1]),
    .b(al_11033702[1]),
    .c(al_42574dc6),
    .o({al_56f6746e,al_c67bebad[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc96c084 (
    .a(al_1315ed94[37]),
    .b(al_11033702[37]),
    .c(al_9a3c1ab7),
    .o({al_16b85269,al_c67bebad[37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc93f476 (
    .a(al_1315ed94[38]),
    .b(al_11033702[38]),
    .c(al_16b85269),
    .o({al_38249694,al_c67bebad[38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bea0d2b8 (
    .a(al_1315ed94[39]),
    .b(al_11033702[39]),
    .c(al_38249694),
    .o({al_f6144b57,al_c67bebad[39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_368990f0 (
    .a(al_1315ed94[40]),
    .b(al_11033702[40]),
    .c(al_f6144b57),
    .o({al_6da3c5cb,al_c67bebad[40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ba912dab (
    .a(al_1315ed94[41]),
    .b(al_11033702[41]),
    .c(al_6da3c5cb),
    .o({al_996323c0,al_c67bebad[41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a081c0b2 (
    .a(al_1315ed94[42]),
    .b(al_11033702[42]),
    .c(al_996323c0),
    .o({al_edd3bfe4,al_c67bebad[42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_458b8f4d (
    .a(al_1315ed94[43]),
    .b(al_11033702[43]),
    .c(al_edd3bfe4),
    .o({al_440c7d0a,al_c67bebad[43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b724ba6 (
    .a(al_1315ed94[44]),
    .b(al_11033702[44]),
    .c(al_440c7d0a),
    .o({al_4629f076,al_c67bebad[44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_64750080 (
    .a(al_1315ed94[45]),
    .b(al_11033702[45]),
    .c(al_4629f076),
    .o({al_689ae363,al_c67bebad[45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_63e240d6 (
    .a(al_1315ed94[46]),
    .b(al_11033702[46]),
    .c(al_689ae363),
    .o({al_d264df46,al_c67bebad[46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_1315ed94[2]),
    .b(al_11033702[2]),
    .c(al_56f6746e),
    .o({al_62cc2266,al_c67bebad[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_39822f5e (
    .a(al_1315ed94[47]),
    .b(al_11033702[47]),
    .c(al_d264df46),
    .o({al_29fe8473,al_c67bebad[47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_298d4cb8 (
    .a(al_1315ed94[48]),
    .b(al_11033702[48]),
    .c(al_29fe8473),
    .o({al_a0aced5d,al_c67bebad[48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_313635c6 (
    .a(al_1315ed94[49]),
    .b(al_11033702[49]),
    .c(al_a0aced5d),
    .o({al_bd3178ec,al_c67bebad[49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_440f6d6d (
    .a(al_1315ed94[50]),
    .b(al_11033702[50]),
    .c(al_bd3178ec),
    .o({al_2a30141f,al_c67bebad[50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef4f93a6 (
    .a(al_1315ed94[51]),
    .b(al_11033702[51]),
    .c(al_2a30141f),
    .o({al_e391dfd4,al_c67bebad[51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8e93da27 (
    .a(al_1315ed94[52]),
    .b(al_11033702[52]),
    .c(al_e391dfd4),
    .o({al_c31d4d4f,al_c67bebad[52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_955595a3 (
    .a(al_1315ed94[53]),
    .b(al_11033702[53]),
    .c(al_c31d4d4f),
    .o({al_432a2e5b,al_c67bebad[53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b31da46b (
    .a(al_1315ed94[54]),
    .b(al_11033702[54]),
    .c(al_432a2e5b),
    .o({al_59ff8a59,al_c67bebad[54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dfd4a7b0 (
    .a(al_1315ed94[55]),
    .b(al_11033702[55]),
    .c(al_59ff8a59),
    .o({al_c27564f1,al_c67bebad[55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a23a824 (
    .a(al_1315ed94[56]),
    .b(al_11033702[56]),
    .c(al_c27564f1),
    .o({al_dcd01a2d,al_c67bebad[56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_1315ed94[3]),
    .b(al_11033702[3]),
    .c(al_62cc2266),
    .o({al_3be447ce,al_c67bebad[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40fca01c (
    .a(al_1315ed94[57]),
    .b(al_11033702[57]),
    .c(al_dcd01a2d),
    .o({al_9d2f5762,al_c67bebad[57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7fc49024 (
    .a(al_1315ed94[58]),
    .b(al_11033702[58]),
    .c(al_9d2f5762),
    .o({al_7cb87941,al_c67bebad[58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce2d27ed (
    .a(al_1315ed94[59]),
    .b(al_11033702[59]),
    .c(al_7cb87941),
    .o({al_5c338988,al_c67bebad[59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e8c29e5 (
    .a(al_1315ed94[60]),
    .b(al_11033702[60]),
    .c(al_5c338988),
    .o({al_9040c841,al_c67bebad[60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8c86c74b (
    .a(al_1315ed94[61]),
    .b(al_11033702[61]),
    .c(al_9040c841),
    .o({al_3f505dba,al_c67bebad[61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b0dd8135 (
    .a(al_1315ed94[62]),
    .b(al_11033702[62]),
    .c(al_3f505dba),
    .o({al_1d0cd6c7,al_c67bebad[62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_22690046 (
    .a(al_1315ed94[63]),
    .b(al_11033702[63]),
    .c(al_1d0cd6c7),
    .o({open_n138,al_c67bebad[63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_1315ed94[4]),
    .b(al_11033702[4]),
    .c(al_3be447ce),
    .o({al_76e76f5,al_c67bebad[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_1315ed94[5]),
    .b(al_11033702[5]),
    .c(al_76e76f5),
    .o({al_40413c0d,al_c67bebad[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_1315ed94[6]),
    .b(al_11033702[6]),
    .c(al_40413c0d),
    .o({al_a2e09ed2,al_c67bebad[6]}));

endmodule 

